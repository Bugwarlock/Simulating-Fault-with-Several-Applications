
//Verilog file of module c6288


`timescale 1 ns / 1ns

module c6288_net(in256,
in239,
in222,
in205,
in188,
in171,
in154,
in137,
in120,
in103,
in86,
in69,
in52,
in35,
in18,
in1,
in528,
in511,
in494,
in477,
in460,
in443,
in426,
in409,
in392,
in375,
in358,
in341,
in324,
in307,
in290,
in273,
out6287,
out6288,
out6280,
out6270,
out6260,
out6250,
out6240,
out6230,
out6220,
out6210,
out6200,
out6190,
out6180,
out6170,
out6160,
out6150,
out6123,
out5971,
out5672,
out5308,
out4946,
out4591,
out4241,
out3895,
out3552,
out3211,
out2877,
out2548,
out2223,
out1901,
out1581,
out545);
  input          in256;
  input          in239;
  input          in222;
  input          in205;
  input          in188;
  input          in171;
  input          in154;
  input          in137;
  input          in120;
  input          in103;
  input          in86;
  input          in69;
  input          in52;
  input          in35;
  input          in18;
  input          in1;
  input          in528;
  input          in511;
  input          in494;
  input          in477;
  input          in460;
  input          in443;
  input          in426;
  input          in409;
  input          in392;
  input          in375;
  input          in358;
  input          in341;
  input          in324;
  input          in307;
  input          in290;
  input          in273;

  output         out6287;
  output         out6288;
  output         out6280;
  output         out6270;
  output         out6260;
  output         out6250;
  output         out6240;
  output         out6230;
  output         out6220;
  output         out6210;
  output         out6200;
  output         out6190;
  output         out6180;
  output         out6170;
  output         out6160;
  output         out6150;
  output         out6123;
  output         out5971;
  output         out5672;
  output         out5308;
  output         out4946;
  output         out4591;
  output         out4241;
  output         out3895;
  output         out3552;
  output         out3211;
  output         out2877;
  output         out2548;
  output         out2223;
  output         out1901;
  output         out1581;
  output         out545;

wire
c6288_wire_1,
c6288_wire_2,
c6288_wire_3,
c6288_wire_4,
c6288_wire_5,
c6288_wire_6,
c6288_wire_7,
c6288_wire_8,
c6288_wire_9,
c6288_wire_10,
c6288_wire_11,
c6288_wire_12,
c6288_wire_13,
c6288_wire_14,
c6288_wire_15,
c6288_wire_16,
c6288_wire_17,
c6288_wire_18,
c6288_wire_19,
c6288_wire_20,
c6288_wire_21,
c6288_wire_22,
c6288_wire_23,
c6288_wire_24,
c6288_wire_25,
c6288_wire_26,
c6288_wire_27,
c6288_wire_28,
c6288_wire_29,
c6288_wire_30,
c6288_wire_31,
c6288_wire_32,
c6288_wire_33,
c6288_wire_34,
c6288_wire_35,
c6288_wire_36,
c6288_wire_37,
c6288_wire_38,
c6288_wire_39,
c6288_wire_40,
c6288_wire_41,
c6288_wire_42,
c6288_wire_43,
c6288_wire_44,
c6288_wire_45,
c6288_wire_46,
c6288_wire_47,
c6288_wire_48,
c6288_wire_49,
c6288_wire_50,
c6288_wire_51,
c6288_wire_52,
c6288_wire_53,
c6288_wire_54,
c6288_wire_55,
c6288_wire_56,
c6288_wire_57,
c6288_wire_58,
c6288_wire_59,
c6288_wire_60,
c6288_wire_61,
c6288_wire_62,
c6288_wire_63,
c6288_wire_64,
c6288_wire_65,
c6288_wire_66,
c6288_wire_67,
c6288_wire_68,
c6288_wire_69,
c6288_wire_70,
c6288_wire_71,
c6288_wire_72,
c6288_wire_73,
c6288_wire_74,
c6288_wire_75,
c6288_wire_76,
c6288_wire_77,
c6288_wire_78,
c6288_wire_79,
c6288_wire_80,
c6288_wire_81,
c6288_wire_82,
c6288_wire_83,
c6288_wire_84,
c6288_wire_85,
c6288_wire_86,
c6288_wire_87,
c6288_wire_88,
c6288_wire_89,
c6288_wire_90,
c6288_wire_91,
c6288_wire_92,
c6288_wire_93,
c6288_wire_94,
c6288_wire_95,
c6288_wire_96,
c6288_wire_97,
c6288_wire_98,
c6288_wire_99,
c6288_wire_100,
c6288_wire_101,
c6288_wire_102,
c6288_wire_103,
c6288_wire_104,
c6288_wire_105,
c6288_wire_106,
c6288_wire_107,
c6288_wire_108,
c6288_wire_109,
c6288_wire_110,
c6288_wire_111,
c6288_wire_112,
c6288_wire_113,
c6288_wire_114,
c6288_wire_115,
c6288_wire_116,
c6288_wire_117,
c6288_wire_118,
c6288_wire_119,
c6288_wire_120,
c6288_wire_121,
c6288_wire_122,
c6288_wire_123,
c6288_wire_124,
c6288_wire_125,
c6288_wire_126,
c6288_wire_127,
c6288_wire_128,
c6288_wire_129,
c6288_wire_130,
c6288_wire_131,
c6288_wire_132,
c6288_wire_133,
c6288_wire_134,
c6288_wire_135,
c6288_wire_136,
c6288_wire_137,
c6288_wire_138,
c6288_wire_139,
c6288_wire_140,
c6288_wire_141,
c6288_wire_142,
c6288_wire_143,
c6288_wire_144,
c6288_wire_145,
c6288_wire_146,
c6288_wire_147,
c6288_wire_148,
c6288_wire_149,
c6288_wire_150,
c6288_wire_151,
c6288_wire_152,
c6288_wire_153,
c6288_wire_154,
c6288_wire_155,
c6288_wire_156,
c6288_wire_157,
c6288_wire_158,
c6288_wire_159,
c6288_wire_160,
c6288_wire_161,
c6288_wire_162,
c6288_wire_163,
c6288_wire_164,
c6288_wire_165,
c6288_wire_166,
c6288_wire_167,
c6288_wire_168,
c6288_wire_169,
c6288_wire_170,
c6288_wire_171,
c6288_wire_172,
c6288_wire_173,
c6288_wire_174,
c6288_wire_175,
c6288_wire_176,
c6288_wire_177,
c6288_wire_178,
c6288_wire_179,
c6288_wire_180,
c6288_wire_181,
c6288_wire_182,
c6288_wire_183,
c6288_wire_184,
c6288_wire_185,
c6288_wire_186,
c6288_wire_187,
c6288_wire_188,
c6288_wire_189,
c6288_wire_190,
c6288_wire_191,
c6288_wire_192,
c6288_wire_193,
c6288_wire_194,
c6288_wire_195,
c6288_wire_196,
c6288_wire_197,
c6288_wire_198,
c6288_wire_199,
c6288_wire_200,
c6288_wire_201,
c6288_wire_202,
c6288_wire_203,
c6288_wire_204,
c6288_wire_205,
c6288_wire_206,
c6288_wire_207,
c6288_wire_208,
c6288_wire_209,
c6288_wire_210,
c6288_wire_211,
c6288_wire_212,
c6288_wire_213,
c6288_wire_214,
c6288_wire_215,
c6288_wire_216,
c6288_wire_217,
c6288_wire_218,
c6288_wire_219,
c6288_wire_220,
c6288_wire_221,
c6288_wire_222,
c6288_wire_223,
c6288_wire_224,
c6288_wire_225,
c6288_wire_226,
c6288_wire_227,
c6288_wire_228,
c6288_wire_229,
c6288_wire_230,
c6288_wire_231,
c6288_wire_232,
c6288_wire_233,
c6288_wire_234,
c6288_wire_235,
c6288_wire_236,
c6288_wire_237,
c6288_wire_238,
c6288_wire_239,
c6288_wire_240,
c6288_wire_241,
c6288_wire_242,
c6288_wire_243,
c6288_wire_244,
c6288_wire_245,
c6288_wire_246,
c6288_wire_247,
c6288_wire_248,
c6288_wire_249,
c6288_wire_250,
c6288_wire_251,
c6288_wire_252,
c6288_wire_253,
c6288_wire_254,
c6288_wire_255,
c6288_wire_256,
c6288_wire_257,
c6288_wire_258,
c6288_wire_259,
c6288_wire_260,
c6288_wire_261,
c6288_wire_262,
c6288_wire_263,
c6288_wire_264,
c6288_wire_265,
c6288_wire_266,
c6288_wire_267,
c6288_wire_268,
c6288_wire_269,
c6288_wire_270,
c6288_wire_271,
c6288_wire_272,
c6288_wire_273,
c6288_wire_274,
c6288_wire_275,
c6288_wire_276,
c6288_wire_277,
c6288_wire_278,
c6288_wire_279,
c6288_wire_280,
c6288_wire_281,
c6288_wire_282,
c6288_wire_283,
c6288_wire_284,
c6288_wire_285,
c6288_wire_286,
c6288_wire_287,
c6288_wire_288,
c6288_wire_289,
c6288_wire_290,
c6288_wire_291,
c6288_wire_292,
c6288_wire_293,
c6288_wire_294,
c6288_wire_295,
c6288_wire_296,
c6288_wire_297,
c6288_wire_298,
c6288_wire_299,
c6288_wire_300,
c6288_wire_301,
c6288_wire_302,
c6288_wire_303,
c6288_wire_304,
c6288_wire_305,
c6288_wire_306,
c6288_wire_307,
c6288_wire_308,
c6288_wire_309,
c6288_wire_310,
c6288_wire_311,
c6288_wire_312,
c6288_wire_313,
c6288_wire_314,
c6288_wire_315,
c6288_wire_316,
c6288_wire_317,
c6288_wire_318,
c6288_wire_319,
c6288_wire_320,
c6288_wire_321,
c6288_wire_322,
c6288_wire_323,
c6288_wire_324,
c6288_wire_325,
c6288_wire_326,
c6288_wire_327,
c6288_wire_328,
c6288_wire_329,
c6288_wire_330,
c6288_wire_331,
c6288_wire_332,
c6288_wire_333,
c6288_wire_334,
c6288_wire_335,
c6288_wire_336,
c6288_wire_337,
c6288_wire_338,
c6288_wire_339,
c6288_wire_340,
c6288_wire_341,
c6288_wire_342,
c6288_wire_343,
c6288_wire_344,
c6288_wire_345,
c6288_wire_346,
c6288_wire_347,
c6288_wire_348,
c6288_wire_349,
c6288_wire_350,
c6288_wire_351,
c6288_wire_352,
c6288_wire_353,
c6288_wire_354,
c6288_wire_355,
c6288_wire_356,
c6288_wire_357,
c6288_wire_358,
c6288_wire_359,
c6288_wire_360,
c6288_wire_361,
c6288_wire_362,
c6288_wire_363,
c6288_wire_364,
c6288_wire_365,
c6288_wire_366,
c6288_wire_367,
c6288_wire_368,
c6288_wire_369,
c6288_wire_370,
c6288_wire_371,
c6288_wire_372,
c6288_wire_373,
c6288_wire_374,
c6288_wire_375,
c6288_wire_376,
c6288_wire_377,
c6288_wire_378,
c6288_wire_379,
c6288_wire_380,
c6288_wire_381,
c6288_wire_382,
c6288_wire_383,
c6288_wire_384,
c6288_wire_385,
c6288_wire_386,
c6288_wire_387,
c6288_wire_388,
c6288_wire_389,
c6288_wire_390,
c6288_wire_391,
c6288_wire_392,
c6288_wire_393,
c6288_wire_394,
c6288_wire_395,
c6288_wire_396,
c6288_wire_397,
c6288_wire_398,
c6288_wire_399,
c6288_wire_400,
c6288_wire_401,
c6288_wire_402,
c6288_wire_403,
c6288_wire_404,
c6288_wire_405,
c6288_wire_406,
c6288_wire_407,
c6288_wire_408,
c6288_wire_409,
c6288_wire_410,
c6288_wire_411,
c6288_wire_412,
c6288_wire_413,
c6288_wire_414,
c6288_wire_415,
c6288_wire_416,
c6288_wire_417,
c6288_wire_418,
c6288_wire_419,
c6288_wire_420,
c6288_wire_421,
c6288_wire_422,
c6288_wire_423,
c6288_wire_424,
c6288_wire_425,
c6288_wire_426,
c6288_wire_427,
c6288_wire_428,
c6288_wire_429,
c6288_wire_430,
c6288_wire_431,
c6288_wire_432,
c6288_wire_433,
c6288_wire_434,
c6288_wire_435,
c6288_wire_436,
c6288_wire_437,
c6288_wire_438,
c6288_wire_439,
c6288_wire_440,
c6288_wire_441,
c6288_wire_442,
c6288_wire_443,
c6288_wire_444,
c6288_wire_445,
c6288_wire_446,
c6288_wire_447,
c6288_wire_448,
c6288_wire_449,
c6288_wire_450,
c6288_wire_451,
c6288_wire_452,
c6288_wire_453,
c6288_wire_454,
c6288_wire_455,
c6288_wire_456,
c6288_wire_457,
c6288_wire_458,
c6288_wire_459,
c6288_wire_460,
c6288_wire_461,
c6288_wire_462,
c6288_wire_463,
c6288_wire_464,
c6288_wire_465,
c6288_wire_466,
c6288_wire_467,
c6288_wire_468,
c6288_wire_469,
c6288_wire_470,
c6288_wire_471,
c6288_wire_472,
c6288_wire_473,
c6288_wire_474,
c6288_wire_475,
c6288_wire_476,
c6288_wire_477,
c6288_wire_478,
c6288_wire_479,
c6288_wire_480,
c6288_wire_481,
c6288_wire_482,
c6288_wire_483,
c6288_wire_484,
c6288_wire_485,
c6288_wire_486,
c6288_wire_487,
c6288_wire_488,
c6288_wire_489,
c6288_wire_490,
c6288_wire_491,
c6288_wire_492,
c6288_wire_493,
c6288_wire_494,
c6288_wire_495,
c6288_wire_496,
c6288_wire_497,
c6288_wire_498,
c6288_wire_499,
c6288_wire_500,
c6288_wire_501,
c6288_wire_502,
c6288_wire_503,
c6288_wire_504,
c6288_wire_505,
c6288_wire_506,
c6288_wire_507,
c6288_wire_508,
c6288_wire_509,
c6288_wire_510,
c6288_wire_511,
c6288_wire_512,
c6288_wire_513,
c6288_wire_514,
c6288_wire_515,
c6288_wire_516,
c6288_wire_517,
c6288_wire_518,
c6288_wire_519,
c6288_wire_520,
c6288_wire_521,
c6288_wire_522,
c6288_wire_523,
c6288_wire_524,
c6288_wire_525,
c6288_wire_526,
c6288_wire_527,
c6288_wire_528,
c6288_wire_529,
c6288_wire_530,
c6288_wire_531,
c6288_wire_532,
c6288_wire_533,
c6288_wire_534,
c6288_wire_535,
c6288_wire_536,
c6288_wire_537,
c6288_wire_538,
c6288_wire_539,
c6288_wire_540,
c6288_wire_541,
c6288_wire_542,
c6288_wire_543,
c6288_wire_544,
c6288_wire_545,
c6288_wire_546,
c6288_wire_547,
c6288_wire_548,
c6288_wire_549,
c6288_wire_550,
c6288_wire_551,
c6288_wire_552,
c6288_wire_553,
c6288_wire_554,
c6288_wire_555,
c6288_wire_556,
c6288_wire_557,
c6288_wire_558,
c6288_wire_559,
c6288_wire_560,
c6288_wire_561,
c6288_wire_562,
c6288_wire_563,
c6288_wire_564,
c6288_wire_565,
c6288_wire_566,
c6288_wire_567,
c6288_wire_568,
c6288_wire_569,
c6288_wire_570,
c6288_wire_571,
c6288_wire_572,
c6288_wire_573,
c6288_wire_574,
c6288_wire_575,
c6288_wire_576,
c6288_wire_577,
c6288_wire_578,
c6288_wire_579,
c6288_wire_580,
c6288_wire_581,
c6288_wire_582,
c6288_wire_583,
c6288_wire_584,
c6288_wire_585,
c6288_wire_586,
c6288_wire_587,
c6288_wire_588,
c6288_wire_589,
c6288_wire_590,
c6288_wire_591,
c6288_wire_592,
c6288_wire_593,
c6288_wire_594,
c6288_wire_595,
c6288_wire_596,
c6288_wire_597,
c6288_wire_598,
c6288_wire_599,
c6288_wire_600,
c6288_wire_601,
c6288_wire_602,
c6288_wire_603,
c6288_wire_604,
c6288_wire_605,
c6288_wire_606,
c6288_wire_607,
c6288_wire_608,
c6288_wire_609,
c6288_wire_610,
c6288_wire_611,
c6288_wire_612,
c6288_wire_613,
c6288_wire_614,
c6288_wire_615,
c6288_wire_616,
c6288_wire_617,
c6288_wire_618,
c6288_wire_619,
c6288_wire_620,
c6288_wire_621,
c6288_wire_622,
c6288_wire_623,
c6288_wire_624,
c6288_wire_625,
c6288_wire_626,
c6288_wire_627,
c6288_wire_628,
c6288_wire_629,
c6288_wire_630,
c6288_wire_631,
c6288_wire_632,
c6288_wire_633,
c6288_wire_634,
c6288_wire_635,
c6288_wire_636,
c6288_wire_637,
c6288_wire_638,
c6288_wire_639,
c6288_wire_640,
c6288_wire_641,
c6288_wire_642,
c6288_wire_643,
c6288_wire_644,
c6288_wire_645,
c6288_wire_646,
c6288_wire_647,
c6288_wire_648,
c6288_wire_649,
c6288_wire_650,
c6288_wire_651,
c6288_wire_652,
c6288_wire_653,
c6288_wire_654,
c6288_wire_655,
c6288_wire_656,
c6288_wire_657,
c6288_wire_658,
c6288_wire_659,
c6288_wire_660,
c6288_wire_661,
c6288_wire_662,
c6288_wire_663,
c6288_wire_664,
c6288_wire_665,
c6288_wire_666,
c6288_wire_667,
c6288_wire_668,
c6288_wire_669,
c6288_wire_670,
c6288_wire_671,
c6288_wire_672,
c6288_wire_673,
c6288_wire_674,
c6288_wire_675,
c6288_wire_676,
c6288_wire_677,
c6288_wire_678,
c6288_wire_679,
c6288_wire_680,
c6288_wire_681,
c6288_wire_682,
c6288_wire_683,
c6288_wire_684,
c6288_wire_685,
c6288_wire_686,
c6288_wire_687,
c6288_wire_688,
c6288_wire_689,
c6288_wire_690,
c6288_wire_691,
c6288_wire_692,
c6288_wire_693,
c6288_wire_694,
c6288_wire_695,
c6288_wire_696,
c6288_wire_697,
c6288_wire_698,
c6288_wire_699,
c6288_wire_700,
c6288_wire_701,
c6288_wire_702,
c6288_wire_703,
c6288_wire_704,
c6288_wire_705,
c6288_wire_706,
c6288_wire_707,
c6288_wire_708,
c6288_wire_709,
c6288_wire_710,
c6288_wire_711,
c6288_wire_712,
c6288_wire_713,
c6288_wire_714,
c6288_wire_715,
c6288_wire_716,
c6288_wire_717,
c6288_wire_718,
c6288_wire_719,
c6288_wire_720,
c6288_wire_721,
c6288_wire_722,
c6288_wire_723,
c6288_wire_724,
c6288_wire_725,
c6288_wire_726,
c6288_wire_727,
c6288_wire_728,
c6288_wire_729,
c6288_wire_730,
c6288_wire_731,
c6288_wire_732,
c6288_wire_733,
c6288_wire_734,
c6288_wire_735,
c6288_wire_736,
c6288_wire_737,
c6288_wire_738,
c6288_wire_739,
c6288_wire_740,
c6288_wire_741,
c6288_wire_742,
c6288_wire_743,
c6288_wire_744,
c6288_wire_745,
c6288_wire_746,
c6288_wire_747,
c6288_wire_748,
c6288_wire_749,
c6288_wire_750,
c6288_wire_751,
c6288_wire_752,
c6288_wire_753,
c6288_wire_754,
c6288_wire_755,
c6288_wire_756,
c6288_wire_757,
c6288_wire_758,
c6288_wire_759,
c6288_wire_760,
c6288_wire_761,
c6288_wire_762,
c6288_wire_763,
c6288_wire_764,
c6288_wire_765,
c6288_wire_766,
c6288_wire_767,
c6288_wire_768,
c6288_wire_769,
c6288_wire_770,
c6288_wire_771,
c6288_wire_772,
c6288_wire_773,
c6288_wire_774,
c6288_wire_775,
c6288_wire_776,
c6288_wire_777,
c6288_wire_778,
c6288_wire_779,
c6288_wire_780,
c6288_wire_781,
c6288_wire_782,
c6288_wire_783,
c6288_wire_784,
c6288_wire_785,
c6288_wire_786,
c6288_wire_787,
c6288_wire_788,
c6288_wire_789,
c6288_wire_790,
c6288_wire_791,
c6288_wire_792,
c6288_wire_793,
c6288_wire_794,
c6288_wire_795,
c6288_wire_796,
c6288_wire_797,
c6288_wire_798,
c6288_wire_799,
c6288_wire_800,
c6288_wire_801,
c6288_wire_802,
c6288_wire_803,
c6288_wire_804,
c6288_wire_805,
c6288_wire_806,
c6288_wire_807,
c6288_wire_808,
c6288_wire_809,
c6288_wire_810,
c6288_wire_811,
c6288_wire_812,
c6288_wire_813,
c6288_wire_814,
c6288_wire_815,
c6288_wire_816,
c6288_wire_817,
c6288_wire_818,
c6288_wire_819,
c6288_wire_820,
c6288_wire_821,
c6288_wire_822,
c6288_wire_823,
c6288_wire_824,
c6288_wire_825,
c6288_wire_826,
c6288_wire_827,
c6288_wire_828,
c6288_wire_829,
c6288_wire_830,
c6288_wire_831,
c6288_wire_832,
c6288_wire_833,
c6288_wire_834,
c6288_wire_835,
c6288_wire_836,
c6288_wire_837,
c6288_wire_838,
c6288_wire_839,
c6288_wire_840,
c6288_wire_841,
c6288_wire_842,
c6288_wire_843,
c6288_wire_844,
c6288_wire_845,
c6288_wire_846,
c6288_wire_847,
c6288_wire_848,
c6288_wire_849,
c6288_wire_850,
c6288_wire_851,
c6288_wire_852,
c6288_wire_853,
c6288_wire_854,
c6288_wire_855,
c6288_wire_856,
c6288_wire_857,
c6288_wire_858,
c6288_wire_859,
c6288_wire_860,
c6288_wire_861,
c6288_wire_862,
c6288_wire_863,
c6288_wire_864,
c6288_wire_865,
c6288_wire_866,
c6288_wire_867,
c6288_wire_868,
c6288_wire_869,
c6288_wire_870,
c6288_wire_871,
c6288_wire_872,
c6288_wire_873,
c6288_wire_874,
c6288_wire_875,
c6288_wire_876,
c6288_wire_877,
c6288_wire_878,
c6288_wire_879,
c6288_wire_880,
c6288_wire_881,
c6288_wire_882,
c6288_wire_883,
c6288_wire_884,
c6288_wire_885,
c6288_wire_886,
c6288_wire_887,
c6288_wire_888,
c6288_wire_889,
c6288_wire_890,
c6288_wire_891,
c6288_wire_892,
c6288_wire_893,
c6288_wire_894,
c6288_wire_895,
c6288_wire_896,
c6288_wire_897,
c6288_wire_898,
c6288_wire_899,
c6288_wire_900,
c6288_wire_901,
c6288_wire_902,
c6288_wire_903,
c6288_wire_904,
c6288_wire_905,
c6288_wire_906,
c6288_wire_907,
c6288_wire_908,
c6288_wire_909,
c6288_wire_910,
c6288_wire_911,
c6288_wire_912,
c6288_wire_913,
c6288_wire_914,
c6288_wire_915,
c6288_wire_916,
c6288_wire_917,
c6288_wire_918,
c6288_wire_919,
c6288_wire_920,
c6288_wire_921,
c6288_wire_922,
c6288_wire_923,
c6288_wire_924,
c6288_wire_925,
c6288_wire_926,
c6288_wire_927,
c6288_wire_928,
c6288_wire_929,
c6288_wire_930,
c6288_wire_931,
c6288_wire_932,
c6288_wire_933,
c6288_wire_934,
c6288_wire_935,
c6288_wire_936,
c6288_wire_937,
c6288_wire_938,
c6288_wire_939,
c6288_wire_940,
c6288_wire_941,
c6288_wire_942,
c6288_wire_943,
c6288_wire_944,
c6288_wire_945,
c6288_wire_946,
c6288_wire_947,
c6288_wire_948,
c6288_wire_949,
c6288_wire_950,
c6288_wire_951,
c6288_wire_952,
c6288_wire_953,
c6288_wire_954,
c6288_wire_955,
c6288_wire_956,
c6288_wire_957,
c6288_wire_958,
c6288_wire_959,
c6288_wire_960,
c6288_wire_961,
c6288_wire_962,
c6288_wire_963,
c6288_wire_964,
c6288_wire_965,
c6288_wire_966,
c6288_wire_967,
c6288_wire_968,
c6288_wire_969,
c6288_wire_970,
c6288_wire_971,
c6288_wire_972,
c6288_wire_973,
c6288_wire_974,
c6288_wire_975,
c6288_wire_976,
c6288_wire_977,
c6288_wire_978,
c6288_wire_979,
c6288_wire_980,
c6288_wire_981,
c6288_wire_982,
c6288_wire_983,
c6288_wire_984,
c6288_wire_985,
c6288_wire_986,
c6288_wire_987,
c6288_wire_988,
c6288_wire_989,
c6288_wire_990,
c6288_wire_991,
c6288_wire_992,
c6288_wire_993,
c6288_wire_994,
c6288_wire_995,
c6288_wire_996,
c6288_wire_997,
c6288_wire_998,
c6288_wire_999,
c6288_wire_1000,
c6288_wire_1001,
c6288_wire_1002,
c6288_wire_1003,
c6288_wire_1004,
c6288_wire_1005,
c6288_wire_1006,
c6288_wire_1007,
c6288_wire_1008,
c6288_wire_1009,
c6288_wire_1010,
c6288_wire_1011,
c6288_wire_1012,
c6288_wire_1013,
c6288_wire_1014,
c6288_wire_1015,
c6288_wire_1016,
c6288_wire_1017,
c6288_wire_1018,
c6288_wire_1019,
c6288_wire_1020,
c6288_wire_1021,
c6288_wire_1022,
c6288_wire_1023,
c6288_wire_1024,
c6288_wire_1025,
c6288_wire_1026,
c6288_wire_1027,
c6288_wire_1028,
c6288_wire_1029,
c6288_wire_1030,
c6288_wire_1031,
c6288_wire_1032,
c6288_wire_1033,
c6288_wire_1034,
c6288_wire_1035,
c6288_wire_1036,
c6288_wire_1037,
c6288_wire_1038,
c6288_wire_1039,
c6288_wire_1040,
c6288_wire_1041,
c6288_wire_1042,
c6288_wire_1043,
c6288_wire_1044,
c6288_wire_1045,
c6288_wire_1046,
c6288_wire_1047,
c6288_wire_1048,
c6288_wire_1049,
c6288_wire_1050,
c6288_wire_1051,
c6288_wire_1052,
c6288_wire_1053,
c6288_wire_1054,
c6288_wire_1055,
c6288_wire_1056,
c6288_wire_1057,
c6288_wire_1058,
c6288_wire_1059,
c6288_wire_1060,
c6288_wire_1061,
c6288_wire_1062,
c6288_wire_1063,
c6288_wire_1064,
c6288_wire_1065,
c6288_wire_1066,
c6288_wire_1067,
c6288_wire_1068,
c6288_wire_1069,
c6288_wire_1070,
c6288_wire_1071,
c6288_wire_1072,
c6288_wire_1073,
c6288_wire_1074,
c6288_wire_1075,
c6288_wire_1076,
c6288_wire_1077,
c6288_wire_1078,
c6288_wire_1079,
c6288_wire_1080,
c6288_wire_1081,
c6288_wire_1082,
c6288_wire_1083,
c6288_wire_1084,
c6288_wire_1085,
c6288_wire_1086,
c6288_wire_1087,
c6288_wire_1088,
c6288_wire_1089,
c6288_wire_1090,
c6288_wire_1091,
c6288_wire_1092,
c6288_wire_1093,
c6288_wire_1094,
c6288_wire_1095,
c6288_wire_1096,
c6288_wire_1097,
c6288_wire_1098,
c6288_wire_1099,
c6288_wire_1100,
c6288_wire_1101,
c6288_wire_1102,
c6288_wire_1103,
c6288_wire_1104,
c6288_wire_1105,
c6288_wire_1106,
c6288_wire_1107,
c6288_wire_1108,
c6288_wire_1109,
c6288_wire_1110,
c6288_wire_1111,
c6288_wire_1112,
c6288_wire_1113,
c6288_wire_1114,
c6288_wire_1115,
c6288_wire_1116,
c6288_wire_1117,
c6288_wire_1118,
c6288_wire_1119,
c6288_wire_1120,
c6288_wire_1121,
c6288_wire_1122,
c6288_wire_1123,
c6288_wire_1124,
c6288_wire_1125,
c6288_wire_1126,
c6288_wire_1127,
c6288_wire_1128,
c6288_wire_1129,
c6288_wire_1130,
c6288_wire_1131,
c6288_wire_1132,
c6288_wire_1133,
c6288_wire_1134,
c6288_wire_1135,
c6288_wire_1136,
c6288_wire_1137,
c6288_wire_1138,
c6288_wire_1139,
c6288_wire_1140,
c6288_wire_1141,
c6288_wire_1142,
c6288_wire_1143,
c6288_wire_1144,
c6288_wire_1145,
c6288_wire_1146,
c6288_wire_1147,
c6288_wire_1148,
c6288_wire_1149,
c6288_wire_1150,
c6288_wire_1151,
c6288_wire_1152,
c6288_wire_1153,
c6288_wire_1154,
c6288_wire_1155,
c6288_wire_1156,
c6288_wire_1157,
c6288_wire_1158,
c6288_wire_1159,
c6288_wire_1160,
c6288_wire_1161,
c6288_wire_1162,
c6288_wire_1163,
c6288_wire_1164,
c6288_wire_1165,
c6288_wire_1166,
c6288_wire_1167,
c6288_wire_1168,
c6288_wire_1169,
c6288_wire_1170,
c6288_wire_1171,
c6288_wire_1172,
c6288_wire_1173,
c6288_wire_1174,
c6288_wire_1175,
c6288_wire_1176,
c6288_wire_1177,
c6288_wire_1178,
c6288_wire_1179,
c6288_wire_1180,
c6288_wire_1181,
c6288_wire_1182,
c6288_wire_1183,
c6288_wire_1184,
c6288_wire_1185,
c6288_wire_1186,
c6288_wire_1187,
c6288_wire_1188,
c6288_wire_1189,
c6288_wire_1190,
c6288_wire_1191,
c6288_wire_1192,
c6288_wire_1193,
c6288_wire_1194,
c6288_wire_1195,
c6288_wire_1196,
c6288_wire_1197,
c6288_wire_1198,
c6288_wire_1199,
c6288_wire_1200,
c6288_wire_1201,
c6288_wire_1202,
c6288_wire_1203,
c6288_wire_1204,
c6288_wire_1205,
c6288_wire_1206,
c6288_wire_1207,
c6288_wire_1208,
c6288_wire_1209,
c6288_wire_1210,
c6288_wire_1211,
c6288_wire_1212,
c6288_wire_1213,
c6288_wire_1214,
c6288_wire_1215,
c6288_wire_1216,
c6288_wire_1217,
c6288_wire_1218,
c6288_wire_1219,
c6288_wire_1220,
c6288_wire_1221,
c6288_wire_1222,
c6288_wire_1223,
c6288_wire_1224,
c6288_wire_1225,
c6288_wire_1226,
c6288_wire_1227,
c6288_wire_1228,
c6288_wire_1229,
c6288_wire_1230,
c6288_wire_1231,
c6288_wire_1232,
c6288_wire_1233,
c6288_wire_1234,
c6288_wire_1235,
c6288_wire_1236,
c6288_wire_1237,
c6288_wire_1238,
c6288_wire_1239,
c6288_wire_1240,
c6288_wire_1241,
c6288_wire_1242,
c6288_wire_1243,
c6288_wire_1244,
c6288_wire_1245,
c6288_wire_1246,
c6288_wire_1247,
c6288_wire_1248,
c6288_wire_1249,
c6288_wire_1250,
c6288_wire_1251,
c6288_wire_1252,
c6288_wire_1253,
c6288_wire_1254,
c6288_wire_1255,
c6288_wire_1256,
c6288_wire_1257,
c6288_wire_1258,
c6288_wire_1259,
c6288_wire_1260,
c6288_wire_1261,
c6288_wire_1262,
c6288_wire_1263,
c6288_wire_1264,
c6288_wire_1265,
c6288_wire_1266,
c6288_wire_1267,
c6288_wire_1268,
c6288_wire_1269,
c6288_wire_1270,
c6288_wire_1271,
c6288_wire_1272,
c6288_wire_1273,
c6288_wire_1274,
c6288_wire_1275,
c6288_wire_1276,
c6288_wire_1277,
c6288_wire_1278,
c6288_wire_1279,
c6288_wire_1280,
c6288_wire_1281,
c6288_wire_1282,
c6288_wire_1283,
c6288_wire_1284,
c6288_wire_1285,
c6288_wire_1286,
c6288_wire_1287,
c6288_wire_1288,
c6288_wire_1289,
c6288_wire_1290,
c6288_wire_1291,
c6288_wire_1292,
c6288_wire_1293,
c6288_wire_1294,
c6288_wire_1295,
c6288_wire_1296,
c6288_wire_1297,
c6288_wire_1298,
c6288_wire_1299,
c6288_wire_1300,
c6288_wire_1301,
c6288_wire_1302,
c6288_wire_1303,
c6288_wire_1304,
c6288_wire_1305,
c6288_wire_1306,
c6288_wire_1307,
c6288_wire_1308,
c6288_wire_1309,
c6288_wire_1310,
c6288_wire_1311,
c6288_wire_1312,
c6288_wire_1313,
c6288_wire_1314,
c6288_wire_1315,
c6288_wire_1316,
c6288_wire_1317,
c6288_wire_1318,
c6288_wire_1319,
c6288_wire_1320,
c6288_wire_1321,
c6288_wire_1322,
c6288_wire_1323,
c6288_wire_1324,
c6288_wire_1325,
c6288_wire_1326,
c6288_wire_1327,
c6288_wire_1328,
c6288_wire_1329,
c6288_wire_1330,
c6288_wire_1331,
c6288_wire_1332,
c6288_wire_1333,
c6288_wire_1334,
c6288_wire_1335,
c6288_wire_1336,
c6288_wire_1337,
c6288_wire_1338,
c6288_wire_1339,
c6288_wire_1340,
c6288_wire_1341,
c6288_wire_1342,
c6288_wire_1343,
c6288_wire_1344,
c6288_wire_1345,
c6288_wire_1346,
c6288_wire_1347,
c6288_wire_1348,
c6288_wire_1349,
c6288_wire_1350,
c6288_wire_1351,
c6288_wire_1352,
c6288_wire_1353,
c6288_wire_1354,
c6288_wire_1355,
c6288_wire_1356,
c6288_wire_1357,
c6288_wire_1358,
c6288_wire_1359,
c6288_wire_1360,
c6288_wire_1361,
c6288_wire_1362,
c6288_wire_1363,
c6288_wire_1364,
c6288_wire_1365,
c6288_wire_1366,
c6288_wire_1367,
c6288_wire_1368,
c6288_wire_1369,
c6288_wire_1370,
c6288_wire_1371,
c6288_wire_1372,
c6288_wire_1373,
c6288_wire_1374,
c6288_wire_1375,
c6288_wire_1376,
c6288_wire_1377,
c6288_wire_1378,
c6288_wire_1379,
c6288_wire_1380,
c6288_wire_1381,
c6288_wire_1382,
c6288_wire_1383,
c6288_wire_1384,
c6288_wire_1385,
c6288_wire_1386,
c6288_wire_1387,
c6288_wire_1388,
c6288_wire_1389,
c6288_wire_1390,
c6288_wire_1391,
c6288_wire_1392,
c6288_wire_1393,
c6288_wire_1394,
c6288_wire_1395,
c6288_wire_1396,
c6288_wire_1397,
c6288_wire_1398,
c6288_wire_1399,
c6288_wire_1400,
c6288_wire_1401,
c6288_wire_1402,
c6288_wire_1403,
c6288_wire_1404,
c6288_wire_1405,
c6288_wire_1406,
c6288_wire_1407,
c6288_wire_1408,
c6288_wire_1409,
c6288_wire_1410,
c6288_wire_1411,
c6288_wire_1412,
c6288_wire_1413,
c6288_wire_1414,
c6288_wire_1415,
c6288_wire_1416,
c6288_wire_1417,
c6288_wire_1418,
c6288_wire_1419,
c6288_wire_1420,
c6288_wire_1421,
c6288_wire_1422,
c6288_wire_1423,
c6288_wire_1424,
c6288_wire_1425,
c6288_wire_1426,
c6288_wire_1427,
c6288_wire_1428,
c6288_wire_1429,
c6288_wire_1430,
c6288_wire_1431,
c6288_wire_1432,
c6288_wire_1433,
c6288_wire_1434,
c6288_wire_1435,
c6288_wire_1436,
c6288_wire_1437,
c6288_wire_1438,
c6288_wire_1439,
c6288_wire_1440,
c6288_wire_1441,
c6288_wire_1442,
c6288_wire_1443,
c6288_wire_1444,
c6288_wire_1445,
c6288_wire_1446,
c6288_wire_1447,
c6288_wire_1448,
c6288_wire_1449,
c6288_wire_1450,
c6288_wire_1451,
c6288_wire_1452,
c6288_wire_1453,
c6288_wire_1454,
c6288_wire_1455,
c6288_wire_1456,
c6288_wire_1457,
c6288_wire_1458,
c6288_wire_1459,
c6288_wire_1460,
c6288_wire_1461,
c6288_wire_1462,
c6288_wire_1463,
c6288_wire_1464,
c6288_wire_1465,
c6288_wire_1466,
c6288_wire_1467,
c6288_wire_1468,
c6288_wire_1469,
c6288_wire_1470,
c6288_wire_1471,
c6288_wire_1472,
c6288_wire_1473,
c6288_wire_1474,
c6288_wire_1475,
c6288_wire_1476,
c6288_wire_1477,
c6288_wire_1478,
c6288_wire_1479,
c6288_wire_1480,
c6288_wire_1481,
c6288_wire_1482,
c6288_wire_1483,
c6288_wire_1484,
c6288_wire_1485,
c6288_wire_1486,
c6288_wire_1487,
c6288_wire_1488,
c6288_wire_1489,
c6288_wire_1490,
c6288_wire_1491,
c6288_wire_1492,
c6288_wire_1493,
c6288_wire_1494,
c6288_wire_1495,
c6288_wire_1496,
c6288_wire_1497,
c6288_wire_1498,
c6288_wire_1499,
c6288_wire_1500,
c6288_wire_1501,
c6288_wire_1502,
c6288_wire_1503,
c6288_wire_1504,
c6288_wire_1505,
c6288_wire_1506,
c6288_wire_1507,
c6288_wire_1508,
c6288_wire_1509,
c6288_wire_1510,
c6288_wire_1511,
c6288_wire_1512,
c6288_wire_1513,
c6288_wire_1514,
c6288_wire_1515,
c6288_wire_1516,
c6288_wire_1517,
c6288_wire_1518,
c6288_wire_1519,
c6288_wire_1520,
c6288_wire_1521,
c6288_wire_1522,
c6288_wire_1523,
c6288_wire_1524,
c6288_wire_1525,
c6288_wire_1526,
c6288_wire_1527,
c6288_wire_1528,
c6288_wire_1529,
c6288_wire_1530,
c6288_wire_1531,
c6288_wire_1532,
c6288_wire_1533,
c6288_wire_1534,
c6288_wire_1535,
c6288_wire_1536,
c6288_wire_1537,
c6288_wire_1538,
c6288_wire_1539,
c6288_wire_1540,
c6288_wire_1541,
c6288_wire_1542,
c6288_wire_1543,
c6288_wire_1544,
c6288_wire_1545,
c6288_wire_1546,
c6288_wire_1547,
c6288_wire_1548,
c6288_wire_1549,
c6288_wire_1550,
c6288_wire_1551,
c6288_wire_1552,
c6288_wire_1553,
c6288_wire_1554,
c6288_wire_1555,
c6288_wire_1556,
c6288_wire_1557,
c6288_wire_1558,
c6288_wire_1559,
c6288_wire_1560,
c6288_wire_1561,
c6288_wire_1562,
c6288_wire_1563,
c6288_wire_1564,
c6288_wire_1565,
c6288_wire_1566,
c6288_wire_1567,
c6288_wire_1568,
c6288_wire_1569,
c6288_wire_1570,
c6288_wire_1571,
c6288_wire_1572,
c6288_wire_1573,
c6288_wire_1574,
c6288_wire_1575,
c6288_wire_1576,
c6288_wire_1577,
c6288_wire_1578,
c6288_wire_1579,
c6288_wire_1580,
c6288_wire_1581,
c6288_wire_1582,
c6288_wire_1583,
c6288_wire_1584,
c6288_wire_1585,
c6288_wire_1586,
c6288_wire_1587,
c6288_wire_1588,
c6288_wire_1589,
c6288_wire_1590,
c6288_wire_1591,
c6288_wire_1592,
c6288_wire_1593,
c6288_wire_1594,
c6288_wire_1595,
c6288_wire_1596,
c6288_wire_1597,
c6288_wire_1598,
c6288_wire_1599,
c6288_wire_1600,
c6288_wire_1601,
c6288_wire_1602,
c6288_wire_1603,
c6288_wire_1604,
c6288_wire_1605,
c6288_wire_1606,
c6288_wire_1607,
c6288_wire_1608,
c6288_wire_1609,
c6288_wire_1610,
c6288_wire_1611,
c6288_wire_1612,
c6288_wire_1613,
c6288_wire_1614,
c6288_wire_1615,
c6288_wire_1616,
c6288_wire_1617,
c6288_wire_1618,
c6288_wire_1619,
c6288_wire_1620,
c6288_wire_1621,
c6288_wire_1622,
c6288_wire_1623,
c6288_wire_1624,
c6288_wire_1625,
c6288_wire_1626,
c6288_wire_1627,
c6288_wire_1628,
c6288_wire_1629,
c6288_wire_1630,
c6288_wire_1631,
c6288_wire_1632,
c6288_wire_1633,
c6288_wire_1634,
c6288_wire_1635,
c6288_wire_1636,
c6288_wire_1637,
c6288_wire_1638,
c6288_wire_1639,
c6288_wire_1640,
c6288_wire_1641,
c6288_wire_1642,
c6288_wire_1643,
c6288_wire_1644,
c6288_wire_1645,
c6288_wire_1646,
c6288_wire_1647,
c6288_wire_1648,
c6288_wire_1649,
c6288_wire_1650,
c6288_wire_1651,
c6288_wire_1652,
c6288_wire_1653,
c6288_wire_1654,
c6288_wire_1655,
c6288_wire_1656,
c6288_wire_1657,
c6288_wire_1658,
c6288_wire_1659,
c6288_wire_1660,
c6288_wire_1661,
c6288_wire_1662,
c6288_wire_1663,
c6288_wire_1664,
c6288_wire_1665,
c6288_wire_1666,
c6288_wire_1667,
c6288_wire_1668,
c6288_wire_1669,
c6288_wire_1670,
c6288_wire_1671,
c6288_wire_1672,
c6288_wire_1673,
c6288_wire_1674,
c6288_wire_1675,
c6288_wire_1676,
c6288_wire_1677,
c6288_wire_1678,
c6288_wire_1679,
c6288_wire_1680,
c6288_wire_1681,
c6288_wire_1682,
c6288_wire_1683,
c6288_wire_1684,
c6288_wire_1685,
c6288_wire_1686,
c6288_wire_1687,
c6288_wire_1688,
c6288_wire_1689,
c6288_wire_1690,
c6288_wire_1691,
c6288_wire_1692,
c6288_wire_1693,
c6288_wire_1694,
c6288_wire_1695,
c6288_wire_1696,
c6288_wire_1697,
c6288_wire_1698,
c6288_wire_1699,
c6288_wire_1700,
c6288_wire_1701,
c6288_wire_1702,
c6288_wire_1703,
c6288_wire_1704,
c6288_wire_1705,
c6288_wire_1706,
c6288_wire_1707,
c6288_wire_1708,
c6288_wire_1709,
c6288_wire_1710,
c6288_wire_1711,
c6288_wire_1712,
c6288_wire_1713,
c6288_wire_1714,
c6288_wire_1715,
c6288_wire_1716,
c6288_wire_1717,
c6288_wire_1718,
c6288_wire_1719,
c6288_wire_1720,
c6288_wire_1721,
c6288_wire_1722,
c6288_wire_1723,
c6288_wire_1724,
c6288_wire_1725,
c6288_wire_1726,
c6288_wire_1727,
c6288_wire_1728,
c6288_wire_1729,
c6288_wire_1730,
c6288_wire_1731,
c6288_wire_1732,
c6288_wire_1733,
c6288_wire_1734,
c6288_wire_1735,
c6288_wire_1736,
c6288_wire_1737,
c6288_wire_1738,
c6288_wire_1739,
c6288_wire_1740,
c6288_wire_1741,
c6288_wire_1742,
c6288_wire_1743,
c6288_wire_1744,
c6288_wire_1745,
c6288_wire_1746,
c6288_wire_1747,
c6288_wire_1748,
c6288_wire_1749,
c6288_wire_1750,
c6288_wire_1751,
c6288_wire_1752,
c6288_wire_1753,
c6288_wire_1754,
c6288_wire_1755,
c6288_wire_1756,
c6288_wire_1757,
c6288_wire_1758,
c6288_wire_1759,
c6288_wire_1760,
c6288_wire_1761,
c6288_wire_1762,
c6288_wire_1763,
c6288_wire_1764,
c6288_wire_1765,
c6288_wire_1766,
c6288_wire_1767,
c6288_wire_1768,
c6288_wire_1769,
c6288_wire_1770,
c6288_wire_1771,
c6288_wire_1772,
c6288_wire_1773,
c6288_wire_1774,
c6288_wire_1775,
c6288_wire_1776,
c6288_wire_1777,
c6288_wire_1778,
c6288_wire_1779,
c6288_wire_1780,
c6288_wire_1781,
c6288_wire_1782,
c6288_wire_1783,
c6288_wire_1784,
c6288_wire_1785,
c6288_wire_1786,
c6288_wire_1787,
c6288_wire_1788,
c6288_wire_1789,
c6288_wire_1790,
c6288_wire_1791,
c6288_wire_1792,
c6288_wire_1793,
c6288_wire_1794,
c6288_wire_1795,
c6288_wire_1796,
c6288_wire_1797,
c6288_wire_1798,
c6288_wire_1799,
c6288_wire_1800,
c6288_wire_1801,
c6288_wire_1802,
c6288_wire_1803,
c6288_wire_1804,
c6288_wire_1805,
c6288_wire_1806,
c6288_wire_1807,
c6288_wire_1808,
c6288_wire_1809,
c6288_wire_1810,
c6288_wire_1811,
c6288_wire_1812,
c6288_wire_1813,
c6288_wire_1814,
c6288_wire_1815,
c6288_wire_1816,
c6288_wire_1817,
c6288_wire_1818,
c6288_wire_1819,
c6288_wire_1820,
c6288_wire_1821,
c6288_wire_1822,
c6288_wire_1823,
c6288_wire_1824,
c6288_wire_1825,
c6288_wire_1826,
c6288_wire_1827,
c6288_wire_1828,
c6288_wire_1829,
c6288_wire_1830,
c6288_wire_1831,
c6288_wire_1832,
c6288_wire_1833,
c6288_wire_1834,
c6288_wire_1835,
c6288_wire_1836,
c6288_wire_1837,
c6288_wire_1838,
c6288_wire_1839,
c6288_wire_1840,
c6288_wire_1841,
c6288_wire_1842,
c6288_wire_1843,
c6288_wire_1844,
c6288_wire_1845,
c6288_wire_1846,
c6288_wire_1847,
c6288_wire_1848,
c6288_wire_1849,
c6288_wire_1850,
c6288_wire_1851,
c6288_wire_1852,
c6288_wire_1853,
c6288_wire_1854,
c6288_wire_1855,
c6288_wire_1856,
c6288_wire_1857,
c6288_wire_1858,
c6288_wire_1859,
c6288_wire_1860,
c6288_wire_1861,
c6288_wire_1862,
c6288_wire_1863,
c6288_wire_1864,
c6288_wire_1865,
c6288_wire_1866,
c6288_wire_1867,
c6288_wire_1868,
c6288_wire_1869,
c6288_wire_1870,
c6288_wire_1871,
c6288_wire_1872,
c6288_wire_1873,
c6288_wire_1874,
c6288_wire_1875,
c6288_wire_1876,
c6288_wire_1877,
c6288_wire_1878,
c6288_wire_1879,
c6288_wire_1880,
c6288_wire_1881,
c6288_wire_1882,
c6288_wire_1883,
c6288_wire_1884,
c6288_wire_1885,
c6288_wire_1886,
c6288_wire_1887,
c6288_wire_1888,
c6288_wire_1889,
c6288_wire_1890,
c6288_wire_1891,
c6288_wire_1892,
c6288_wire_1893,
c6288_wire_1894,
c6288_wire_1895,
c6288_wire_1896,
c6288_wire_1897,
c6288_wire_1898,
c6288_wire_1899,
c6288_wire_1900,
c6288_wire_1901,
c6288_wire_1902,
c6288_wire_1903,
c6288_wire_1904,
c6288_wire_1905,
c6288_wire_1906,
c6288_wire_1907,
c6288_wire_1908,
c6288_wire_1909,
c6288_wire_1910,
c6288_wire_1911,
c6288_wire_1912,
c6288_wire_1913,
c6288_wire_1914,
c6288_wire_1915,
c6288_wire_1916,
c6288_wire_1917,
c6288_wire_1918,
c6288_wire_1919,
c6288_wire_1920,
c6288_wire_1921,
c6288_wire_1922,
c6288_wire_1923,
c6288_wire_1924,
c6288_wire_1925,
c6288_wire_1926,
c6288_wire_1927,
c6288_wire_1928,
c6288_wire_1929,
c6288_wire_1930,
c6288_wire_1931,
c6288_wire_1932,
c6288_wire_1933,
c6288_wire_1934,
c6288_wire_1935,
c6288_wire_1936,
c6288_wire_1937,
c6288_wire_1938,
c6288_wire_1939,
c6288_wire_1940,
c6288_wire_1941,
c6288_wire_1942,
c6288_wire_1943,
c6288_wire_1944,
c6288_wire_1945,
c6288_wire_1946,
c6288_wire_1947,
c6288_wire_1948,
c6288_wire_1949,
c6288_wire_1950,
c6288_wire_1951,
c6288_wire_1952,
c6288_wire_1953,
c6288_wire_1954,
c6288_wire_1955,
c6288_wire_1956,
c6288_wire_1957,
c6288_wire_1958,
c6288_wire_1959,
c6288_wire_1960,
c6288_wire_1961,
c6288_wire_1962,
c6288_wire_1963,
c6288_wire_1964,
c6288_wire_1965,
c6288_wire_1966,
c6288_wire_1967,
c6288_wire_1968,
c6288_wire_1969,
c6288_wire_1970,
c6288_wire_1971,
c6288_wire_1972,
c6288_wire_1973,
c6288_wire_1974,
c6288_wire_1975,
c6288_wire_1976,
c6288_wire_1977,
c6288_wire_1978,
c6288_wire_1979,
c6288_wire_1980,
c6288_wire_1981,
c6288_wire_1982,
c6288_wire_1983,
c6288_wire_1984,
c6288_wire_1985,
c6288_wire_1986,
c6288_wire_1987,
c6288_wire_1988,
c6288_wire_1989,
c6288_wire_1990,
c6288_wire_1991,
c6288_wire_1992,
c6288_wire_1993,
c6288_wire_1994,
c6288_wire_1995,
c6288_wire_1996,
c6288_wire_1997,
c6288_wire_1998,
c6288_wire_1999,
c6288_wire_2000,
c6288_wire_2001,
c6288_wire_2002,
c6288_wire_2003,
c6288_wire_2004,
c6288_wire_2005,
c6288_wire_2006,
c6288_wire_2007,
c6288_wire_2008,
c6288_wire_2009,
c6288_wire_2010,
c6288_wire_2011,
c6288_wire_2012,
c6288_wire_2013,
c6288_wire_2014,
c6288_wire_2015,
c6288_wire_2016,
c6288_wire_2017,
c6288_wire_2018,
c6288_wire_2019,
c6288_wire_2020,
c6288_wire_2021,
c6288_wire_2022,
c6288_wire_2023,
c6288_wire_2024,
c6288_wire_2025,
c6288_wire_2026,
c6288_wire_2027,
c6288_wire_2028,
c6288_wire_2029,
c6288_wire_2030,
c6288_wire_2031,
c6288_wire_2032,
c6288_wire_2033,
c6288_wire_2034,
c6288_wire_2035,
c6288_wire_2036,
c6288_wire_2037,
c6288_wire_2038,
c6288_wire_2039,
c6288_wire_2040,
c6288_wire_2041,
c6288_wire_2042,
c6288_wire_2043,
c6288_wire_2044,
c6288_wire_2045,
c6288_wire_2046,
c6288_wire_2047,
c6288_wire_2048,
c6288_wire_2049,
c6288_wire_2050,
c6288_wire_2051,
c6288_wire_2052,
c6288_wire_2053,
c6288_wire_2054,
c6288_wire_2055,
c6288_wire_2056,
c6288_wire_2057,
c6288_wire_2058,
c6288_wire_2059,
c6288_wire_2060,
c6288_wire_2061,
c6288_wire_2062,
c6288_wire_2063,
c6288_wire_2064,
c6288_wire_2065,
c6288_wire_2066,
c6288_wire_2067,
c6288_wire_2068,
c6288_wire_2069,
c6288_wire_2070,
c6288_wire_2071,
c6288_wire_2072,
c6288_wire_2073,
c6288_wire_2074,
c6288_wire_2075,
c6288_wire_2076,
c6288_wire_2077,
c6288_wire_2078,
c6288_wire_2079,
c6288_wire_2080,
c6288_wire_2081,
c6288_wire_2082,
c6288_wire_2083,
c6288_wire_2084,
c6288_wire_2085,
c6288_wire_2086,
c6288_wire_2087,
c6288_wire_2088,
c6288_wire_2089,
c6288_wire_2090,
c6288_wire_2091,
c6288_wire_2092,
c6288_wire_2093,
c6288_wire_2094,
c6288_wire_2095,
c6288_wire_2096,
c6288_wire_2097,
c6288_wire_2098,
c6288_wire_2099,
c6288_wire_2100,
c6288_wire_2101,
c6288_wire_2102,
c6288_wire_2103,
c6288_wire_2104,
c6288_wire_2105,
c6288_wire_2106,
c6288_wire_2107,
c6288_wire_2108,
c6288_wire_2109,
c6288_wire_2110,
c6288_wire_2111,
c6288_wire_2112,
c6288_wire_2113,
c6288_wire_2114,
c6288_wire_2115,
c6288_wire_2116,
c6288_wire_2117,
c6288_wire_2118,
c6288_wire_2119,
c6288_wire_2120,
c6288_wire_2121,
c6288_wire_2122,
c6288_wire_2123,
c6288_wire_2124,
c6288_wire_2125,
c6288_wire_2126,
c6288_wire_2127,
c6288_wire_2128,
c6288_wire_2129,
c6288_wire_2130,
c6288_wire_2131,
c6288_wire_2132,
c6288_wire_2133,
c6288_wire_2134,
c6288_wire_2135,
c6288_wire_2136,
c6288_wire_2137,
c6288_wire_2138,
c6288_wire_2139,
c6288_wire_2140,
c6288_wire_2141,
c6288_wire_2142,
c6288_wire_2143,
c6288_wire_2144,
c6288_wire_2145,
c6288_wire_2146,
c6288_wire_2147,
c6288_wire_2148,
c6288_wire_2149,
c6288_wire_2150,
c6288_wire_2151,
c6288_wire_2152,
c6288_wire_2153,
c6288_wire_2154,
c6288_wire_2155,
c6288_wire_2156,
c6288_wire_2157,
c6288_wire_2158,
c6288_wire_2159,
c6288_wire_2160,
c6288_wire_2161,
c6288_wire_2162,
c6288_wire_2163,
c6288_wire_2164,
c6288_wire_2165,
c6288_wire_2166,
c6288_wire_2167,
c6288_wire_2168,
c6288_wire_2169,
c6288_wire_2170,
c6288_wire_2171,
c6288_wire_2172,
c6288_wire_2173,
c6288_wire_2174,
c6288_wire_2175,
c6288_wire_2176,
c6288_wire_2177,
c6288_wire_2178,
c6288_wire_2179,
c6288_wire_2180,
c6288_wire_2181,
c6288_wire_2182,
c6288_wire_2183,
c6288_wire_2184,
c6288_wire_2185,
c6288_wire_2186,
c6288_wire_2187,
c6288_wire_2188,
c6288_wire_2189,
c6288_wire_2190,
c6288_wire_2191,
c6288_wire_2192,
c6288_wire_2193,
c6288_wire_2194,
c6288_wire_2195,
c6288_wire_2196,
c6288_wire_2197,
c6288_wire_2198,
c6288_wire_2199,
c6288_wire_2200,
c6288_wire_2201,
c6288_wire_2202,
c6288_wire_2203,
c6288_wire_2204,
c6288_wire_2205,
c6288_wire_2206,
c6288_wire_2207,
c6288_wire_2208,
c6288_wire_2209,
c6288_wire_2210,
c6288_wire_2211,
c6288_wire_2212,
c6288_wire_2213,
c6288_wire_2214,
c6288_wire_2215,
c6288_wire_2216,
c6288_wire_2217,
c6288_wire_2218,
c6288_wire_2219,
c6288_wire_2220,
c6288_wire_2221,
c6288_wire_2222,
c6288_wire_2223,
c6288_wire_2224,
c6288_wire_2225,
c6288_wire_2226,
c6288_wire_2227,
c6288_wire_2228,
c6288_wire_2229,
c6288_wire_2230,
c6288_wire_2231,
c6288_wire_2232,
c6288_wire_2233,
c6288_wire_2234,
c6288_wire_2235,
c6288_wire_2236,
c6288_wire_2237,
c6288_wire_2238,
c6288_wire_2239,
c6288_wire_2240,
c6288_wire_2241,
c6288_wire_2242,
c6288_wire_2243,
c6288_wire_2244,
c6288_wire_2245,
c6288_wire_2246,
c6288_wire_2247,
c6288_wire_2248,
c6288_wire_2249,
c6288_wire_2250,
c6288_wire_2251,
c6288_wire_2252,
c6288_wire_2253,
c6288_wire_2254,
c6288_wire_2255,
c6288_wire_2256,
c6288_wire_2257,
c6288_wire_2258,
c6288_wire_2259,
c6288_wire_2260,
c6288_wire_2261,
c6288_wire_2262,
c6288_wire_2263,
c6288_wire_2264,
c6288_wire_2265,
c6288_wire_2266,
c6288_wire_2267,
c6288_wire_2268,
c6288_wire_2269,
c6288_wire_2270,
c6288_wire_2271,
c6288_wire_2272,
c6288_wire_2273,
c6288_wire_2274,
c6288_wire_2275,
c6288_wire_2276,
c6288_wire_2277,
c6288_wire_2278,
c6288_wire_2279,
c6288_wire_2280,
c6288_wire_2281,
c6288_wire_2282,
c6288_wire_2283,
c6288_wire_2284,
c6288_wire_2285,
c6288_wire_2286,
c6288_wire_2287,
c6288_wire_2288,
c6288_wire_2289,
c6288_wire_2290,
c6288_wire_2291,
c6288_wire_2292,
c6288_wire_2293,
c6288_wire_2294,
c6288_wire_2295,
c6288_wire_2296,
c6288_wire_2297,
c6288_wire_2298,
c6288_wire_2299,
c6288_wire_2300,
c6288_wire_2301,
c6288_wire_2302,
c6288_wire_2303,
c6288_wire_2304,
c6288_wire_2305,
c6288_wire_2306,
c6288_wire_2307,
c6288_wire_2308,
c6288_wire_2309,
c6288_wire_2310,
c6288_wire_2311,
c6288_wire_2312,
c6288_wire_2313,
c6288_wire_2314,
c6288_wire_2315,
c6288_wire_2316,
c6288_wire_2317,
c6288_wire_2318,
c6288_wire_2319,
c6288_wire_2320,
c6288_wire_2321,
c6288_wire_2322,
c6288_wire_2323,
c6288_wire_2324,
c6288_wire_2325,
c6288_wire_2326,
c6288_wire_2327,
c6288_wire_2328,
c6288_wire_2329,
c6288_wire_2330,
c6288_wire_2331,
c6288_wire_2332,
c6288_wire_2333,
c6288_wire_2334,
c6288_wire_2335,
c6288_wire_2336,
c6288_wire_2337,
c6288_wire_2338,
c6288_wire_2339,
c6288_wire_2340,
c6288_wire_2341,
c6288_wire_2342,
c6288_wire_2343,
c6288_wire_2344,
c6288_wire_2345,
c6288_wire_2346,
c6288_wire_2347,
c6288_wire_2348,
c6288_wire_2349,
c6288_wire_2350,
c6288_wire_2351,
c6288_wire_2352,
c6288_wire_2353,
c6288_wire_2354,
c6288_wire_2355,
c6288_wire_2356,
c6288_wire_2357,
c6288_wire_2358,
c6288_wire_2359,
c6288_wire_2360,
c6288_wire_2361,
c6288_wire_2362,
c6288_wire_2363,
c6288_wire_2364,
c6288_wire_2365,
c6288_wire_2366,
c6288_wire_2367,
c6288_wire_2368,
c6288_wire_2369,
c6288_wire_2370,
c6288_wire_2371,
c6288_wire_2372,
c6288_wire_2373,
c6288_wire_2374,
c6288_wire_2375,
c6288_wire_2376,
c6288_wire_2377,
c6288_wire_2378,
c6288_wire_2379,
c6288_wire_2380,
c6288_wire_2381,
c6288_wire_2382,
c6288_wire_2383,
c6288_wire_2384,
c6288_wire_2385,
c6288_wire_2386,
c6288_wire_2387,
c6288_wire_2388,
c6288_wire_2389,
c6288_wire_2390,
c6288_wire_2391,
c6288_wire_2392,
c6288_wire_2393,
c6288_wire_2394,
c6288_wire_2395,
c6288_wire_2396,
c6288_wire_2397,
c6288_wire_2398,
c6288_wire_2399,
c6288_wire_2400,
c6288_wire_2401,
c6288_wire_2402,
c6288_wire_2403,
c6288_wire_2404,
c6288_wire_2405,
c6288_wire_2406,
c6288_wire_2407,
c6288_wire_2408,
c6288_wire_2409,
c6288_wire_2410,
c6288_wire_2411,
c6288_wire_2412,
c6288_wire_2413,
c6288_wire_2414,
c6288_wire_2415,
c6288_wire_2416,
c6288_wire_2417,
c6288_wire_2418,
c6288_wire_2419,
c6288_wire_2420,
c6288_wire_2421,
c6288_wire_2422,
c6288_wire_2423,
c6288_wire_2424,
c6288_wire_2425,
c6288_wire_2426,
c6288_wire_2427,
c6288_wire_2428,
c6288_wire_2429,
c6288_wire_2430,
c6288_wire_2431,
c6288_wire_2432,
c6288_wire_2433,
c6288_wire_2434,
c6288_wire_2435,
c6288_wire_2436,
c6288_wire_2437,
c6288_wire_2438,
c6288_wire_2439,
c6288_wire_2440,
c6288_wire_2441,
c6288_wire_2442,
c6288_wire_2443,
c6288_wire_2444,
c6288_wire_2445,
c6288_wire_2446,
c6288_wire_2447,
c6288_wire_2448,
c6288_wire_2449,
c6288_wire_2450,
c6288_wire_2451,
c6288_wire_2452,
c6288_wire_2453,
c6288_wire_2454,
c6288_wire_2455,
c6288_wire_2456,
c6288_wire_2457,
c6288_wire_2458,
c6288_wire_2459,
c6288_wire_2460,
c6288_wire_2461,
c6288_wire_2462,
c6288_wire_2463,
c6288_wire_2464,
c6288_wire_2465,
c6288_wire_2466,
c6288_wire_2467,
c6288_wire_2468,
c6288_wire_2469,
c6288_wire_2470,
c6288_wire_2471,
c6288_wire_2472,
c6288_wire_2473,
c6288_wire_2474,
c6288_wire_2475,
c6288_wire_2476,
c6288_wire_2477,
c6288_wire_2478,
c6288_wire_2479,
c6288_wire_2480,
c6288_wire_2481,
c6288_wire_2482,
c6288_wire_2483,
c6288_wire_2484,
c6288_wire_2485,
c6288_wire_2486,
c6288_wire_2487,
c6288_wire_2488,
c6288_wire_2489,
c6288_wire_2490,
c6288_wire_2491,
c6288_wire_2492,
c6288_wire_2493,
c6288_wire_2494,
c6288_wire_2495,
c6288_wire_2496,
c6288_wire_2497,
c6288_wire_2498,
c6288_wire_2499,
c6288_wire_2500,
c6288_wire_2501,
c6288_wire_2502,
c6288_wire_2503,
c6288_wire_2504,
c6288_wire_2505,
c6288_wire_2506,
c6288_wire_2507,
c6288_wire_2508,
c6288_wire_2509,
c6288_wire_2510,
c6288_wire_2511,
c6288_wire_2512,
c6288_wire_2513,
c6288_wire_2514,
c6288_wire_2515,
c6288_wire_2516,
c6288_wire_2517,
c6288_wire_2518,
c6288_wire_2519,
c6288_wire_2520,
c6288_wire_2521,
c6288_wire_2522,
c6288_wire_2523,
c6288_wire_2524,
c6288_wire_2525,
c6288_wire_2526,
c6288_wire_2527,
c6288_wire_2528,
c6288_wire_2529,
c6288_wire_2530,
c6288_wire_2531,
c6288_wire_2532,
c6288_wire_2533,
c6288_wire_2534,
c6288_wire_2535,
c6288_wire_2536,
c6288_wire_2537,
c6288_wire_2538,
c6288_wire_2539,
c6288_wire_2540,
c6288_wire_2541,
c6288_wire_2542,
c6288_wire_2543,
c6288_wire_2544,
c6288_wire_2545,
c6288_wire_2546,
c6288_wire_2547,
c6288_wire_2548,
c6288_wire_2549,
c6288_wire_2550,
c6288_wire_2551,
c6288_wire_2552,
c6288_wire_2553,
c6288_wire_2554,
c6288_wire_2555,
c6288_wire_2556,
c6288_wire_2557,
c6288_wire_2558,
c6288_wire_2559,
c6288_wire_2560,
c6288_wire_2561,
c6288_wire_2562,
c6288_wire_2563,
c6288_wire_2564,
c6288_wire_2565,
c6288_wire_2566,
c6288_wire_2567,
c6288_wire_2568,
c6288_wire_2569,
c6288_wire_2570,
c6288_wire_2571,
c6288_wire_2572,
c6288_wire_2573,
c6288_wire_2574,
c6288_wire_2575,
c6288_wire_2576,
c6288_wire_2577,
c6288_wire_2578,
c6288_wire_2579,
c6288_wire_2580,
c6288_wire_2581,
c6288_wire_2582,
c6288_wire_2583,
c6288_wire_2584,
c6288_wire_2585,
c6288_wire_2586,
c6288_wire_2587,
c6288_wire_2588,
c6288_wire_2589,
c6288_wire_2590,
c6288_wire_2591,
c6288_wire_2592,
c6288_wire_2593,
c6288_wire_2594,
c6288_wire_2595,
c6288_wire_2596,
c6288_wire_2597,
c6288_wire_2598,
c6288_wire_2599,
c6288_wire_2600,
c6288_wire_2601,
c6288_wire_2602,
c6288_wire_2603,
c6288_wire_2604,
c6288_wire_2605,
c6288_wire_2606,
c6288_wire_2607,
c6288_wire_2608,
c6288_wire_2609,
c6288_wire_2610,
c6288_wire_2611,
c6288_wire_2612,
c6288_wire_2613,
c6288_wire_2614,
c6288_wire_2615,
c6288_wire_2616,
c6288_wire_2617,
c6288_wire_2618,
c6288_wire_2619,
c6288_wire_2620,
c6288_wire_2621,
c6288_wire_2622,
c6288_wire_2623,
c6288_wire_2624,
c6288_wire_2625,
c6288_wire_2626,
c6288_wire_2627,
c6288_wire_2628,
c6288_wire_2629,
c6288_wire_2630,
c6288_wire_2631,
c6288_wire_2632,
c6288_wire_2633,
c6288_wire_2634,
c6288_wire_2635,
c6288_wire_2636,
c6288_wire_2637,
c6288_wire_2638,
c6288_wire_2639,
c6288_wire_2640,
c6288_wire_2641,
c6288_wire_2642,
c6288_wire_2643,
c6288_wire_2644,
c6288_wire_2645,
c6288_wire_2646,
c6288_wire_2647,
c6288_wire_2648,
c6288_wire_2649,
c6288_wire_2650,
c6288_wire_2651,
c6288_wire_2652,
c6288_wire_2653,
c6288_wire_2654,
c6288_wire_2655,
c6288_wire_2656,
c6288_wire_2657,
c6288_wire_2658,
c6288_wire_2659,
c6288_wire_2660,
c6288_wire_2661,
c6288_wire_2662,
c6288_wire_2663,
c6288_wire_2664,
c6288_wire_2665,
c6288_wire_2666,
c6288_wire_2667,
c6288_wire_2668,
c6288_wire_2669,
c6288_wire_2670,
c6288_wire_2671,
c6288_wire_2672,
c6288_wire_2673,
c6288_wire_2674,
c6288_wire_2675,
c6288_wire_2676,
c6288_wire_2677,
c6288_wire_2678,
c6288_wire_2679,
c6288_wire_2680,
c6288_wire_2681,
c6288_wire_2682,
c6288_wire_2683,
c6288_wire_2684,
c6288_wire_2685,
c6288_wire_2686,
c6288_wire_2687,
c6288_wire_2688,
c6288_wire_2689,
c6288_wire_2690,
c6288_wire_2691,
c6288_wire_2692,
c6288_wire_2693,
c6288_wire_2694,
c6288_wire_2695,
c6288_wire_2696,
c6288_wire_2697,
c6288_wire_2698,
c6288_wire_2699,
c6288_wire_2700,
c6288_wire_2701,
c6288_wire_2702,
c6288_wire_2703,
c6288_wire_2704,
c6288_wire_2705,
c6288_wire_2706,
c6288_wire_2707,
c6288_wire_2708,
c6288_wire_2709,
c6288_wire_2710,
c6288_wire_2711,
c6288_wire_2712,
c6288_wire_2713,
c6288_wire_2714,
c6288_wire_2715,
c6288_wire_2716,
c6288_wire_2717,
c6288_wire_2718,
c6288_wire_2719,
c6288_wire_2720,
c6288_wire_2721,
c6288_wire_2722,
c6288_wire_2723,
c6288_wire_2724,
c6288_wire_2725,
c6288_wire_2726,
c6288_wire_2727,
c6288_wire_2728,
c6288_wire_2729,
c6288_wire_2730,
c6288_wire_2731,
c6288_wire_2732,
c6288_wire_2733,
c6288_wire_2734,
c6288_wire_2735,
c6288_wire_2736,
c6288_wire_2737,
c6288_wire_2738,
c6288_wire_2739,
c6288_wire_2740,
c6288_wire_2741,
c6288_wire_2742,
c6288_wire_2743,
c6288_wire_2744,
c6288_wire_2745,
c6288_wire_2746,
c6288_wire_2747,
c6288_wire_2748,
c6288_wire_2749,
c6288_wire_2750,
c6288_wire_2751,
c6288_wire_2752,
c6288_wire_2753,
c6288_wire_2754,
c6288_wire_2755,
c6288_wire_2756,
c6288_wire_2757,
c6288_wire_2758,
c6288_wire_2759,
c6288_wire_2760,
c6288_wire_2761,
c6288_wire_2762,
c6288_wire_2763,
c6288_wire_2764,
c6288_wire_2765,
c6288_wire_2766,
c6288_wire_2767,
c6288_wire_2768,
c6288_wire_2769,
c6288_wire_2770,
c6288_wire_2771,
c6288_wire_2772,
c6288_wire_2773,
c6288_wire_2774,
c6288_wire_2775,
c6288_wire_2776,
c6288_wire_2777,
c6288_wire_2778,
c6288_wire_2779,
c6288_wire_2780,
c6288_wire_2781,
c6288_wire_2782,
c6288_wire_2783,
c6288_wire_2784,
c6288_wire_2785,
c6288_wire_2786,
c6288_wire_2787,
c6288_wire_2788,
c6288_wire_2789,
c6288_wire_2790,
c6288_wire_2791,
c6288_wire_2792,
c6288_wire_2793,
c6288_wire_2794,
c6288_wire_2795,
c6288_wire_2796,
c6288_wire_2797,
c6288_wire_2798,
c6288_wire_2799,
c6288_wire_2800,
c6288_wire_2801,
c6288_wire_2802,
c6288_wire_2803,
c6288_wire_2804,
c6288_wire_2805,
c6288_wire_2806,
c6288_wire_2807,
c6288_wire_2808,
c6288_wire_2809,
c6288_wire_2810,
c6288_wire_2811,
c6288_wire_2812,
c6288_wire_2813,
c6288_wire_2814,
c6288_wire_2815,
c6288_wire_2816,
c6288_wire_2817,
c6288_wire_2818,
c6288_wire_2819,
c6288_wire_2820,
c6288_wire_2821,
c6288_wire_2822,
c6288_wire_2823,
c6288_wire_2824,
c6288_wire_2825,
c6288_wire_2826,
c6288_wire_2827,
c6288_wire_2828,
c6288_wire_2829,
c6288_wire_2830,
c6288_wire_2831,
c6288_wire_2832,
c6288_wire_2833,
c6288_wire_2834,
c6288_wire_2835,
c6288_wire_2836,
c6288_wire_2837,
c6288_wire_2838,
c6288_wire_2839,
c6288_wire_2840,
c6288_wire_2841,
c6288_wire_2842,
c6288_wire_2843,
c6288_wire_2844,
c6288_wire_2845,
c6288_wire_2846,
c6288_wire_2847,
c6288_wire_2848,
c6288_wire_2849,
c6288_wire_2850,
c6288_wire_2851,
c6288_wire_2852,
c6288_wire_2853,
c6288_wire_2854,
c6288_wire_2855,
c6288_wire_2856,
c6288_wire_2857,
c6288_wire_2858,
c6288_wire_2859,
c6288_wire_2860,
c6288_wire_2861,
c6288_wire_2862,
c6288_wire_2863,
c6288_wire_2864,
c6288_wire_2865,
c6288_wire_2866,
c6288_wire_2867,
c6288_wire_2868,
c6288_wire_2869,
c6288_wire_2870,
c6288_wire_2871,
c6288_wire_2872,
c6288_wire_2873,
c6288_wire_2874,
c6288_wire_2875,
c6288_wire_2876,
c6288_wire_2877,
c6288_wire_2878,
c6288_wire_2879,
c6288_wire_2880,
c6288_wire_2881,
c6288_wire_2882,
c6288_wire_2883,
c6288_wire_2884,
c6288_wire_2885,
c6288_wire_2886,
c6288_wire_2887,
c6288_wire_2888,
c6288_wire_2889,
c6288_wire_2890,
c6288_wire_1_0,
c6288_wire_1_1,
c6288_wire_1_2,
c6288_wire_4_0,
c6288_wire_4_1,
c6288_wire_4_2,
c6288_wire_9_0,
c6288_wire_9_1,
c6288_wire_9_2,
c6288_wire_11_0,
c6288_wire_11_1,
c6288_wire_11_2,
c6288_wire_14_0,
c6288_wire_14_1,
c6288_wire_14_2,
c6288_wire_16_0,
c6288_wire_16_1,
c6288_wire_16_2,
c6288_wire_19_0,
c6288_wire_19_1,
c6288_wire_19_2,
c6288_wire_21_0,
c6288_wire_21_1,
c6288_wire_21_2,
c6288_wire_24_0,
c6288_wire_24_1,
c6288_wire_24_2,
c6288_wire_26_0,
c6288_wire_26_1,
c6288_wire_29_0,
c6288_wire_29_1,
c6288_wire_29_2,
c6288_wire_31_0,
c6288_wire_31_1,
c6288_wire_31_2,
c6288_wire_36_0,
c6288_wire_36_1,
c6288_wire_36_2,
c6288_wire_38_0,
c6288_wire_38_1,
c6288_wire_38_2,
c6288_wire_41_0,
c6288_wire_41_1,
c6288_wire_41_2,
c6288_wire_43_0,
c6288_wire_43_1,
c6288_wire_43_2,
c6288_wire_46_0,
c6288_wire_46_1,
c6288_wire_46_2,
c6288_wire_48_0,
c6288_wire_48_1,
c6288_wire_48_2,
c6288_wire_51_0,
c6288_wire_51_1,
c6288_wire_51_2,
c6288_wire_53_0,
c6288_wire_53_1,
c6288_wire_53_2,
c6288_wire_56_0,
c6288_wire_56_1,
c6288_wire_56_2,
c6288_wire_58_0,
c6288_wire_58_1,
c6288_wire_58_2,
c6288_wire_61_0,
c6288_wire_61_1,
c6288_wire_61_2,
c6288_wire_63_0,
c6288_wire_63_1,
c6288_wire_63_2,
c6288_wire_66_0,
c6288_wire_66_1,
c6288_wire_66_2,
c6288_wire_68_0,
c6288_wire_68_1,
c6288_wire_68_2,
c6288_wire_71_0,
c6288_wire_71_1,
c6288_wire_71_2,
c6288_wire_72_0,
c6288_wire_72_1,
c6288_wire_72_2,
c6288_wire_327_0,
c6288_wire_327_1,
c6288_wire_327_2,
c6288_wire_748_0,
c6288_wire_748_1,
c6288_wire_748_2,
c6288_wire_749_0,
c6288_wire_749_1,
c6288_wire_757_0,
c6288_wire_757_1,
c6288_wire_757_2,
c6288_wire_758_0,
c6288_wire_758_1,
c6288_wire_763_0,
c6288_wire_763_1,
c6288_wire_763_2,
c6288_wire_764_0,
c6288_wire_764_1,
c6288_wire_769_0,
c6288_wire_769_1,
c6288_wire_769_2,
c6288_wire_770_0,
c6288_wire_770_1,
c6288_wire_776_0,
c6288_wire_776_1,
c6288_wire_780_0,
c6288_wire_780_1,
c6288_wire_784_0,
c6288_wire_784_1,
c6288_wire_784_2,
c6288_wire_785_0,
c6288_wire_785_1,
c6288_wire_791_0,
c6288_wire_791_1,
c6288_wire_791_2,
c6288_wire_792_0,
c6288_wire_792_1,
c6288_wire_797_0,
c6288_wire_797_1,
c6288_wire_797_2,
c6288_wire_798_0,
c6288_wire_798_1,
c6288_wire_803_0,
c6288_wire_803_1,
c6288_wire_803_2,
c6288_wire_804_0,
c6288_wire_804_1,
c6288_wire_809_0,
c6288_wire_809_1,
c6288_wire_809_2,
c6288_wire_810_0,
c6288_wire_810_1,
c6288_wire_815_0,
c6288_wire_815_1,
c6288_wire_815_2,
c6288_wire_816_0,
c6288_wire_816_1,
c6288_wire_821_0,
c6288_wire_821_1,
c6288_wire_821_2,
c6288_wire_822_0,
c6288_wire_822_1,
c6288_wire_827_0,
c6288_wire_827_1,
c6288_wire_827_2,
c6288_wire_828_0,
c6288_wire_828_1,
c6288_wire_833_0,
c6288_wire_833_1,
c6288_wire_833_2,
c6288_wire_754_0,
c6288_wire_754_1,
c6288_wire_140_0,
c6288_wire_140_1,
c6288_wire_140_2,
c6288_wire_839_0,
c6288_wire_839_1,
c6288_wire_138_0,
c6288_wire_138_1,
c6288_wire_138_2,
c6288_wire_847_0,
c6288_wire_847_1,
c6288_wire_136_0,
c6288_wire_136_1,
c6288_wire_136_2,
c6288_wire_852_0,
c6288_wire_852_1,
c6288_wire_134_0,
c6288_wire_134_1,
c6288_wire_134_2,
c6288_wire_857_0,
c6288_wire_857_1,
c6288_wire_862_0,
c6288_wire_862_1,
c6288_wire_862_2,
c6288_wire_863_0,
c6288_wire_863_1,
c6288_wire_869_0,
c6288_wire_869_1,
c6288_wire_869_2,
c6288_wire_158_0,
c6288_wire_158_1,
c6288_wire_158_2,
c6288_wire_874_0,
c6288_wire_874_1,
c6288_wire_156_0,
c6288_wire_156_1,
c6288_wire_156_2,
c6288_wire_880_0,
c6288_wire_880_1,
c6288_wire_154_0,
c6288_wire_154_1,
c6288_wire_154_2,
c6288_wire_885_0,
c6288_wire_885_1,
c6288_wire_152_0,
c6288_wire_152_1,
c6288_wire_152_2,
c6288_wire_890_0,
c6288_wire_890_1,
c6288_wire_150_0,
c6288_wire_150_1,
c6288_wire_150_2,
c6288_wire_895_0,
c6288_wire_895_1,
c6288_wire_148_0,
c6288_wire_148_1,
c6288_wire_148_2,
c6288_wire_900_0,
c6288_wire_900_1,
c6288_wire_146_0,
c6288_wire_146_1,
c6288_wire_146_2,
c6288_wire_905_0,
c6288_wire_905_1,
c6288_wire_144_0,
c6288_wire_144_1,
c6288_wire_144_2,
c6288_wire_910_0,
c6288_wire_910_1,
c6288_wire_142_0,
c6288_wire_142_1,
c6288_wire_142_2,
c6288_wire_844_0,
c6288_wire_844_1,
c6288_wire_182_0,
c6288_wire_182_1,
c6288_wire_182_2,
c6288_wire_920_0,
c6288_wire_920_1,
c6288_wire_180_0,
c6288_wire_180_1,
c6288_wire_180_2,
c6288_wire_928_0,
c6288_wire_928_1,
c6288_wire_178_0,
c6288_wire_178_1,
c6288_wire_178_2,
c6288_wire_933_0,
c6288_wire_933_1,
c6288_wire_176_0,
c6288_wire_176_1,
c6288_wire_176_2,
c6288_wire_938_0,
c6288_wire_938_1,
c6288_wire_870_0,
c6288_wire_870_1,
c6288_wire_870_2,
c6288_wire_943_0,
c6288_wire_943_1,
c6288_wire_949_0,
c6288_wire_949_1,
c6288_wire_949_2,
c6288_wire_200_0,
c6288_wire_200_1,
c6288_wire_200_2,
c6288_wire_952_0,
c6288_wire_952_1,
c6288_wire_198_0,
c6288_wire_198_1,
c6288_wire_198_2,
c6288_wire_958_0,
c6288_wire_958_1,
c6288_wire_196_0,
c6288_wire_196_1,
c6288_wire_196_2,
c6288_wire_963_0,
c6288_wire_963_1,
c6288_wire_194_0,
c6288_wire_194_1,
c6288_wire_194_2,
c6288_wire_968_0,
c6288_wire_968_1,
c6288_wire_192_0,
c6288_wire_192_1,
c6288_wire_192_2,
c6288_wire_973_0,
c6288_wire_973_1,
c6288_wire_190_0,
c6288_wire_190_1,
c6288_wire_190_2,
c6288_wire_978_0,
c6288_wire_978_1,
c6288_wire_188_0,
c6288_wire_188_1,
c6288_wire_188_2,
c6288_wire_983_0,
c6288_wire_983_1,
c6288_wire_186_0,
c6288_wire_186_1,
c6288_wire_186_2,
c6288_wire_988_0,
c6288_wire_988_1,
c6288_wire_184_0,
c6288_wire_184_1,
c6288_wire_184_2,
c6288_wire_925_0,
c6288_wire_925_1,
c6288_wire_224_0,
c6288_wire_224_1,
c6288_wire_224_2,
c6288_wire_998_0,
c6288_wire_998_1,
c6288_wire_222_0,
c6288_wire_222_1,
c6288_wire_222_2,
c6288_wire_1006_0,
c6288_wire_1006_1,
c6288_wire_220_0,
c6288_wire_220_1,
c6288_wire_220_2,
c6288_wire_1011_0,
c6288_wire_1011_1,
c6288_wire_218_0,
c6288_wire_218_1,
c6288_wire_218_2,
c6288_wire_1016_0,
c6288_wire_1016_1,
c6288_wire_950_0,
c6288_wire_950_1,
c6288_wire_950_2,
c6288_wire_1021_0,
c6288_wire_1021_1,
c6288_wire_1027_0,
c6288_wire_1027_1,
c6288_wire_1027_2,
c6288_wire_242_0,
c6288_wire_242_1,
c6288_wire_242_2,
c6288_wire_1030_0,
c6288_wire_1030_1,
c6288_wire_240_0,
c6288_wire_240_1,
c6288_wire_240_2,
c6288_wire_1036_0,
c6288_wire_1036_1,
c6288_wire_238_0,
c6288_wire_238_1,
c6288_wire_238_2,
c6288_wire_1041_0,
c6288_wire_1041_1,
c6288_wire_236_0,
c6288_wire_236_1,
c6288_wire_236_2,
c6288_wire_1046_0,
c6288_wire_1046_1,
c6288_wire_234_0,
c6288_wire_234_1,
c6288_wire_234_2,
c6288_wire_1051_0,
c6288_wire_1051_1,
c6288_wire_232_0,
c6288_wire_232_1,
c6288_wire_232_2,
c6288_wire_1056_0,
c6288_wire_1056_1,
c6288_wire_230_0,
c6288_wire_230_1,
c6288_wire_230_2,
c6288_wire_1061_0,
c6288_wire_1061_1,
c6288_wire_228_0,
c6288_wire_228_1,
c6288_wire_228_2,
c6288_wire_1066_0,
c6288_wire_1066_1,
c6288_wire_226_0,
c6288_wire_226_1,
c6288_wire_226_2,
c6288_wire_1003_0,
c6288_wire_1003_1,
c6288_wire_286_0,
c6288_wire_286_1,
c6288_wire_286_2,
c6288_wire_266_0,
c6288_wire_266_1,
c6288_wire_266_2,
c6288_wire_1074_0,
c6288_wire_1074_1,
c6288_wire_264_0,
c6288_wire_264_1,
c6288_wire_264_2,
c6288_wire_1082_0,
c6288_wire_1082_1,
c6288_wire_262_0,
c6288_wire_262_1,
c6288_wire_262_2,
c6288_wire_1087_0,
c6288_wire_1087_1,
c6288_wire_260_0,
c6288_wire_260_1,
c6288_wire_260_2,
c6288_wire_1092_0,
c6288_wire_1092_1,
c6288_wire_1028_0,
c6288_wire_1028_1,
c6288_wire_1028_2,
c6288_wire_1097_0,
c6288_wire_1097_1,
c6288_wire_1103_0,
c6288_wire_1103_1,
c6288_wire_1103_2,
c6288_wire_1103_3,
c6288_wire_1108_0,
c6288_wire_1108_1,
c6288_wire_1108_2,
c6288_wire_282_0,
c6288_wire_282_1,
c6288_wire_282_2,
c6288_wire_1115_0,
c6288_wire_1115_1,
c6288_wire_280_0,
c6288_wire_280_1,
c6288_wire_280_2,
c6288_wire_1120_0,
c6288_wire_1120_1,
c6288_wire_278_0,
c6288_wire_278_1,
c6288_wire_278_2,
c6288_wire_1125_0,
c6288_wire_1125_1,
c6288_wire_276_0,
c6288_wire_276_1,
c6288_wire_276_2,
c6288_wire_1130_0,
c6288_wire_1130_1,
c6288_wire_274_0,
c6288_wire_274_1,
c6288_wire_274_2,
c6288_wire_1135_0,
c6288_wire_1135_1,
c6288_wire_272_0,
c6288_wire_272_1,
c6288_wire_272_2,
c6288_wire_1140_0,
c6288_wire_1140_1,
c6288_wire_270_0,
c6288_wire_270_1,
c6288_wire_270_2,
c6288_wire_1145_0,
c6288_wire_1145_1,
c6288_wire_268_0,
c6288_wire_268_1,
c6288_wire_268_2,
c6288_wire_1079_0,
c6288_wire_1079_1,
c6288_wire_1152_0,
c6288_wire_1152_1,
c6288_wire_1152_2,
c6288_wire_1159_0,
c6288_wire_1159_1,
c6288_wire_1159_2,
c6288_wire_1165_0,
c6288_wire_1165_1,
c6288_wire_1165_2,
c6288_wire_1171_0,
c6288_wire_1171_1,
c6288_wire_1171_2,
c6288_wire_1177_0,
c6288_wire_1177_1,
c6288_wire_1177_2,
c6288_wire_1177_3,
c6288_wire_1186_0,
c6288_wire_1186_1,
c6288_wire_1186_2,
c6288_wire_1192_0,
c6288_wire_1192_1,
c6288_wire_1192_2,
c6288_wire_1198_0,
c6288_wire_1198_1,
c6288_wire_1198_2,
c6288_wire_1204_0,
c6288_wire_1204_1,
c6288_wire_1204_2,
c6288_wire_1210_0,
c6288_wire_1210_1,
c6288_wire_1210_2,
c6288_wire_1216_0,
c6288_wire_1216_1,
c6288_wire_1216_2,
c6288_wire_1222_0,
c6288_wire_1222_1,
c6288_wire_1222_2,
c6288_wire_1228_0,
c6288_wire_1228_1,
c6288_wire_1228_2,
c6288_wire_382_0,
c6288_wire_382_1,
c6288_wire_382_2,
c6288_wire_1236_0,
c6288_wire_1236_1,
c6288_wire_380_0,
c6288_wire_380_1,
c6288_wire_380_2,
c6288_wire_1244_0,
c6288_wire_1244_1,
c6288_wire_378_0,
c6288_wire_378_1,
c6288_wire_378_2,
c6288_wire_1249_0,
c6288_wire_1249_1,
c6288_wire_376_0,
c6288_wire_376_1,
c6288_wire_376_2,
c6288_wire_1254_0,
c6288_wire_1254_1,
c6288_wire_782_0,
c6288_wire_782_1,
c6288_wire_1259_0,
c6288_wire_1259_1,
c6288_wire_1265_0,
c6288_wire_1265_1,
c6288_wire_1265_2,
c6288_wire_400_0,
c6288_wire_400_1,
c6288_wire_400_2,
c6288_wire_1269_0,
c6288_wire_1269_1,
c6288_wire_398_0,
c6288_wire_398_1,
c6288_wire_398_2,
c6288_wire_1275_0,
c6288_wire_1275_1,
c6288_wire_396_0,
c6288_wire_396_1,
c6288_wire_396_2,
c6288_wire_1280_0,
c6288_wire_1280_1,
c6288_wire_394_0,
c6288_wire_394_1,
c6288_wire_394_2,
c6288_wire_1285_0,
c6288_wire_1285_1,
c6288_wire_392_0,
c6288_wire_392_1,
c6288_wire_392_2,
c6288_wire_1290_0,
c6288_wire_1290_1,
c6288_wire_390_0,
c6288_wire_390_1,
c6288_wire_390_2,
c6288_wire_1295_0,
c6288_wire_1295_1,
c6288_wire_388_0,
c6288_wire_388_1,
c6288_wire_388_2,
c6288_wire_1300_0,
c6288_wire_1300_1,
c6288_wire_386_0,
c6288_wire_386_1,
c6288_wire_386_2,
c6288_wire_1305_0,
c6288_wire_1305_1,
c6288_wire_384_0,
c6288_wire_384_1,
c6288_wire_384_2,
c6288_wire_1241_0,
c6288_wire_1241_1,
c6288_wire_424_0,
c6288_wire_424_1,
c6288_wire_424_2,
c6288_wire_1315_0,
c6288_wire_1315_1,
c6288_wire_422_0,
c6288_wire_422_1,
c6288_wire_422_2,
c6288_wire_1323_0,
c6288_wire_1323_1,
c6288_wire_420_0,
c6288_wire_420_1,
c6288_wire_420_2,
c6288_wire_1328_0,
c6288_wire_1328_1,
c6288_wire_418_0,
c6288_wire_418_1,
c6288_wire_418_2,
c6288_wire_1333_0,
c6288_wire_1333_1,
c6288_wire_1266_0,
c6288_wire_1266_1,
c6288_wire_1266_2,
c6288_wire_1338_0,
c6288_wire_1338_1,
c6288_wire_1344_0,
c6288_wire_1344_1,
c6288_wire_1344_2,
c6288_wire_442_0,
c6288_wire_442_1,
c6288_wire_442_2,
c6288_wire_1347_0,
c6288_wire_1347_1,
c6288_wire_440_0,
c6288_wire_440_1,
c6288_wire_440_2,
c6288_wire_1353_0,
c6288_wire_1353_1,
c6288_wire_438_0,
c6288_wire_438_1,
c6288_wire_438_2,
c6288_wire_1358_0,
c6288_wire_1358_1,
c6288_wire_436_0,
c6288_wire_436_1,
c6288_wire_436_2,
c6288_wire_1363_0,
c6288_wire_1363_1,
c6288_wire_434_0,
c6288_wire_434_1,
c6288_wire_434_2,
c6288_wire_1368_0,
c6288_wire_1368_1,
c6288_wire_432_0,
c6288_wire_432_1,
c6288_wire_432_2,
c6288_wire_1373_0,
c6288_wire_1373_1,
c6288_wire_430_0,
c6288_wire_430_1,
c6288_wire_430_2,
c6288_wire_1378_0,
c6288_wire_1378_1,
c6288_wire_428_0,
c6288_wire_428_1,
c6288_wire_428_2,
c6288_wire_1383_0,
c6288_wire_1383_1,
c6288_wire_426_0,
c6288_wire_426_1,
c6288_wire_426_2,
c6288_wire_1320_0,
c6288_wire_1320_1,
c6288_wire_466_0,
c6288_wire_466_1,
c6288_wire_466_2,
c6288_wire_1393_0,
c6288_wire_1393_1,
c6288_wire_464_0,
c6288_wire_464_1,
c6288_wire_464_2,
c6288_wire_1401_0,
c6288_wire_1401_1,
c6288_wire_462_0,
c6288_wire_462_1,
c6288_wire_462_2,
c6288_wire_1406_0,
c6288_wire_1406_1,
c6288_wire_460_0,
c6288_wire_460_1,
c6288_wire_460_2,
c6288_wire_1411_0,
c6288_wire_1411_1,
c6288_wire_1345_0,
c6288_wire_1345_1,
c6288_wire_1345_2,
c6288_wire_1416_0,
c6288_wire_1416_1,
c6288_wire_1422_0,
c6288_wire_1422_1,
c6288_wire_1422_2,
c6288_wire_484_0,
c6288_wire_484_1,
c6288_wire_484_2,
c6288_wire_1425_0,
c6288_wire_1425_1,
c6288_wire_482_0,
c6288_wire_482_1,
c6288_wire_482_2,
c6288_wire_1431_0,
c6288_wire_1431_1,
c6288_wire_480_0,
c6288_wire_480_1,
c6288_wire_480_2,
c6288_wire_1436_0,
c6288_wire_1436_1,
c6288_wire_478_0,
c6288_wire_478_1,
c6288_wire_478_2,
c6288_wire_1441_0,
c6288_wire_1441_1,
c6288_wire_476_0,
c6288_wire_476_1,
c6288_wire_476_2,
c6288_wire_1446_0,
c6288_wire_1446_1,
c6288_wire_474_0,
c6288_wire_474_1,
c6288_wire_474_2,
c6288_wire_1451_0,
c6288_wire_1451_1,
c6288_wire_472_0,
c6288_wire_472_1,
c6288_wire_472_2,
c6288_wire_1456_0,
c6288_wire_1456_1,
c6288_wire_470_0,
c6288_wire_470_1,
c6288_wire_470_2,
c6288_wire_1461_0,
c6288_wire_1461_1,
c6288_wire_468_0,
c6288_wire_468_1,
c6288_wire_468_2,
c6288_wire_1398_0,
c6288_wire_1398_1,
c6288_wire_508_0,
c6288_wire_508_1,
c6288_wire_508_2,
c6288_wire_1471_0,
c6288_wire_1471_1,
c6288_wire_506_0,
c6288_wire_506_1,
c6288_wire_506_2,
c6288_wire_1479_0,
c6288_wire_1479_1,
c6288_wire_504_0,
c6288_wire_504_1,
c6288_wire_504_2,
c6288_wire_1484_0,
c6288_wire_1484_1,
c6288_wire_502_0,
c6288_wire_502_1,
c6288_wire_502_2,
c6288_wire_1489_0,
c6288_wire_1489_1,
c6288_wire_1423_0,
c6288_wire_1423_1,
c6288_wire_1423_2,
c6288_wire_1494_0,
c6288_wire_1494_1,
c6288_wire_1500_0,
c6288_wire_1500_1,
c6288_wire_1500_2,
c6288_wire_526_0,
c6288_wire_526_1,
c6288_wire_526_2,
c6288_wire_1503_0,
c6288_wire_1503_1,
c6288_wire_524_0,
c6288_wire_524_1,
c6288_wire_524_2,
c6288_wire_1509_0,
c6288_wire_1509_1,
c6288_wire_522_0,
c6288_wire_522_1,
c6288_wire_522_2,
c6288_wire_1514_0,
c6288_wire_1514_1,
c6288_wire_520_0,
c6288_wire_520_1,
c6288_wire_520_2,
c6288_wire_1519_0,
c6288_wire_1519_1,
c6288_wire_518_0,
c6288_wire_518_1,
c6288_wire_518_2,
c6288_wire_1524_0,
c6288_wire_1524_1,
c6288_wire_516_0,
c6288_wire_516_1,
c6288_wire_516_2,
c6288_wire_1529_0,
c6288_wire_1529_1,
c6288_wire_514_0,
c6288_wire_514_1,
c6288_wire_514_2,
c6288_wire_1534_0,
c6288_wire_1534_1,
c6288_wire_512_0,
c6288_wire_512_1,
c6288_wire_512_2,
c6288_wire_1539_0,
c6288_wire_1539_1,
c6288_wire_510_0,
c6288_wire_510_1,
c6288_wire_510_2,
c6288_wire_1476_0,
c6288_wire_1476_1,
c6288_wire_550_0,
c6288_wire_550_1,
c6288_wire_550_2,
c6288_wire_1549_0,
c6288_wire_1549_1,
c6288_wire_548_0,
c6288_wire_548_1,
c6288_wire_548_2,
c6288_wire_1557_0,
c6288_wire_1557_1,
c6288_wire_546_0,
c6288_wire_546_1,
c6288_wire_546_2,
c6288_wire_1562_0,
c6288_wire_1562_1,
c6288_wire_544_0,
c6288_wire_544_1,
c6288_wire_544_2,
c6288_wire_1567_0,
c6288_wire_1567_1,
c6288_wire_1501_0,
c6288_wire_1501_1,
c6288_wire_1501_2,
c6288_wire_1572_0,
c6288_wire_1572_1,
c6288_wire_1578_0,
c6288_wire_1578_1,
c6288_wire_1578_2,
c6288_wire_568_0,
c6288_wire_568_1,
c6288_wire_568_2,
c6288_wire_1581_0,
c6288_wire_1581_1,
c6288_wire_566_0,
c6288_wire_566_1,
c6288_wire_566_2,
c6288_wire_1587_0,
c6288_wire_1587_1,
c6288_wire_564_0,
c6288_wire_564_1,
c6288_wire_564_2,
c6288_wire_1592_0,
c6288_wire_1592_1,
c6288_wire_562_0,
c6288_wire_562_1,
c6288_wire_562_2,
c6288_wire_1597_0,
c6288_wire_1597_1,
c6288_wire_560_0,
c6288_wire_560_1,
c6288_wire_560_2,
c6288_wire_1602_0,
c6288_wire_1602_1,
c6288_wire_558_0,
c6288_wire_558_1,
c6288_wire_558_2,
c6288_wire_1607_0,
c6288_wire_1607_1,
c6288_wire_556_0,
c6288_wire_556_1,
c6288_wire_556_2,
c6288_wire_1612_0,
c6288_wire_1612_1,
c6288_wire_554_0,
c6288_wire_554_1,
c6288_wire_554_2,
c6288_wire_1617_0,
c6288_wire_1617_1,
c6288_wire_552_0,
c6288_wire_552_1,
c6288_wire_552_2,
c6288_wire_1554_0,
c6288_wire_1554_1,
c6288_wire_592_0,
c6288_wire_592_1,
c6288_wire_592_2,
c6288_wire_1627_0,
c6288_wire_1627_1,
c6288_wire_590_0,
c6288_wire_590_1,
c6288_wire_590_2,
c6288_wire_1635_0,
c6288_wire_1635_1,
c6288_wire_588_0,
c6288_wire_588_1,
c6288_wire_588_2,
c6288_wire_1640_0,
c6288_wire_1640_1,
c6288_wire_586_0,
c6288_wire_586_1,
c6288_wire_586_2,
c6288_wire_1645_0,
c6288_wire_1645_1,
c6288_wire_1579_0,
c6288_wire_1579_1,
c6288_wire_1579_2,
c6288_wire_1650_0,
c6288_wire_1650_1,
c6288_wire_1656_0,
c6288_wire_1656_1,
c6288_wire_1656_2,
c6288_wire_610_0,
c6288_wire_610_1,
c6288_wire_610_2,
c6288_wire_1659_0,
c6288_wire_1659_1,
c6288_wire_608_0,
c6288_wire_608_1,
c6288_wire_608_2,
c6288_wire_1665_0,
c6288_wire_1665_1,
c6288_wire_606_0,
c6288_wire_606_1,
c6288_wire_606_2,
c6288_wire_1670_0,
c6288_wire_1670_1,
c6288_wire_604_0,
c6288_wire_604_1,
c6288_wire_604_2,
c6288_wire_1675_0,
c6288_wire_1675_1,
c6288_wire_602_0,
c6288_wire_602_1,
c6288_wire_602_2,
c6288_wire_1680_0,
c6288_wire_1680_1,
c6288_wire_600_0,
c6288_wire_600_1,
c6288_wire_600_2,
c6288_wire_1685_0,
c6288_wire_1685_1,
c6288_wire_598_0,
c6288_wire_598_1,
c6288_wire_598_2,
c6288_wire_1690_0,
c6288_wire_1690_1,
c6288_wire_596_0,
c6288_wire_596_1,
c6288_wire_596_2,
c6288_wire_1695_0,
c6288_wire_1695_1,
c6288_wire_594_0,
c6288_wire_594_1,
c6288_wire_594_2,
c6288_wire_1632_0,
c6288_wire_1632_1,
c6288_wire_634_0,
c6288_wire_634_1,
c6288_wire_634_2,
c6288_wire_1705_0,
c6288_wire_1705_1,
c6288_wire_632_0,
c6288_wire_632_1,
c6288_wire_632_2,
c6288_wire_1713_0,
c6288_wire_1713_1,
c6288_wire_630_0,
c6288_wire_630_1,
c6288_wire_630_2,
c6288_wire_1718_0,
c6288_wire_1718_1,
c6288_wire_628_0,
c6288_wire_628_1,
c6288_wire_628_2,
c6288_wire_1723_0,
c6288_wire_1723_1,
c6288_wire_1657_0,
c6288_wire_1657_1,
c6288_wire_1657_2,
c6288_wire_1728_0,
c6288_wire_1728_1,
c6288_wire_1734_0,
c6288_wire_1734_1,
c6288_wire_1734_2,
c6288_wire_652_0,
c6288_wire_652_1,
c6288_wire_652_2,
c6288_wire_1737_0,
c6288_wire_1737_1,
c6288_wire_650_0,
c6288_wire_650_1,
c6288_wire_650_2,
c6288_wire_1743_0,
c6288_wire_1743_1,
c6288_wire_648_0,
c6288_wire_648_1,
c6288_wire_648_2,
c6288_wire_1748_0,
c6288_wire_1748_1,
c6288_wire_646_0,
c6288_wire_646_1,
c6288_wire_646_2,
c6288_wire_1753_0,
c6288_wire_1753_1,
c6288_wire_644_0,
c6288_wire_644_1,
c6288_wire_644_2,
c6288_wire_1758_0,
c6288_wire_1758_1,
c6288_wire_642_0,
c6288_wire_642_1,
c6288_wire_642_2,
c6288_wire_1763_0,
c6288_wire_1763_1,
c6288_wire_640_0,
c6288_wire_640_1,
c6288_wire_640_2,
c6288_wire_1768_0,
c6288_wire_1768_1,
c6288_wire_638_0,
c6288_wire_638_1,
c6288_wire_638_2,
c6288_wire_1773_0,
c6288_wire_1773_1,
c6288_wire_636_0,
c6288_wire_636_1,
c6288_wire_636_2,
c6288_wire_1710_0,
c6288_wire_1710_1,
c6288_wire_676_0,
c6288_wire_676_1,
c6288_wire_676_2,
c6288_wire_1783_0,
c6288_wire_1783_1,
c6288_wire_674_0,
c6288_wire_674_1,
c6288_wire_674_2,
c6288_wire_1791_0,
c6288_wire_1791_1,
c6288_wire_672_0,
c6288_wire_672_1,
c6288_wire_672_2,
c6288_wire_1796_0,
c6288_wire_1796_1,
c6288_wire_670_0,
c6288_wire_670_1,
c6288_wire_670_2,
c6288_wire_1801_0,
c6288_wire_1801_1,
c6288_wire_1735_0,
c6288_wire_1735_1,
c6288_wire_1735_2,
c6288_wire_1806_0,
c6288_wire_1806_1,
c6288_wire_1812_0,
c6288_wire_1812_1,
c6288_wire_1812_2,
c6288_wire_694_0,
c6288_wire_694_1,
c6288_wire_694_2,
c6288_wire_1815_0,
c6288_wire_1815_1,
c6288_wire_692_0,
c6288_wire_692_1,
c6288_wire_692_2,
c6288_wire_1821_0,
c6288_wire_1821_1,
c6288_wire_690_0,
c6288_wire_690_1,
c6288_wire_690_2,
c6288_wire_1826_0,
c6288_wire_1826_1,
c6288_wire_688_0,
c6288_wire_688_1,
c6288_wire_688_2,
c6288_wire_1831_0,
c6288_wire_1831_1,
c6288_wire_686_0,
c6288_wire_686_1,
c6288_wire_686_2,
c6288_wire_1836_0,
c6288_wire_1836_1,
c6288_wire_684_0,
c6288_wire_684_1,
c6288_wire_684_2,
c6288_wire_1841_0,
c6288_wire_1841_1,
c6288_wire_682_0,
c6288_wire_682_1,
c6288_wire_682_2,
c6288_wire_1846_0,
c6288_wire_1846_1,
c6288_wire_680_0,
c6288_wire_680_1,
c6288_wire_680_2,
c6288_wire_1851_0,
c6288_wire_1851_1,
c6288_wire_678_0,
c6288_wire_678_1,
c6288_wire_678_2,
c6288_wire_1788_0,
c6288_wire_1788_1,
c6288_wire_718_0,
c6288_wire_718_1,
c6288_wire_718_2,
c6288_wire_1861_0,
c6288_wire_1861_1,
c6288_wire_716_0,
c6288_wire_716_1,
c6288_wire_716_2,
c6288_wire_1869_0,
c6288_wire_1869_1,
c6288_wire_714_0,
c6288_wire_714_1,
c6288_wire_714_2,
c6288_wire_1874_0,
c6288_wire_1874_1,
c6288_wire_712_0,
c6288_wire_712_1,
c6288_wire_712_2,
c6288_wire_1879_0,
c6288_wire_1879_1,
c6288_wire_1813_0,
c6288_wire_1813_1,
c6288_wire_1813_2,
c6288_wire_1884_0,
c6288_wire_1884_1,
c6288_wire_873_0,
c6288_wire_873_1,
c6288_wire_873_2,
c6288_wire_736_0,
c6288_wire_736_1,
c6288_wire_736_2,
c6288_wire_1890_0,
c6288_wire_1890_1,
c6288_wire_734_0,
c6288_wire_734_1,
c6288_wire_734_2,
c6288_wire_1896_0,
c6288_wire_1896_1,
c6288_wire_732_0,
c6288_wire_732_1,
c6288_wire_732_2,
c6288_wire_1901_0,
c6288_wire_1901_1,
c6288_wire_730_0,
c6288_wire_730_1,
c6288_wire_730_2,
c6288_wire_1906_0,
c6288_wire_1906_1,
c6288_wire_728_0,
c6288_wire_728_1,
c6288_wire_728_2,
c6288_wire_1911_0,
c6288_wire_1911_1,
c6288_wire_726_0,
c6288_wire_726_1,
c6288_wire_726_2,
c6288_wire_1916_0,
c6288_wire_1916_1,
c6288_wire_724_0,
c6288_wire_724_1,
c6288_wire_724_2,
c6288_wire_1921_0,
c6288_wire_1921_1,
c6288_wire_722_0,
c6288_wire_722_1,
c6288_wire_722_2,
c6288_wire_1926_0,
c6288_wire_1926_1,
c6288_wire_720_0,
c6288_wire_720_1,
c6288_wire_720_2,
c6288_wire_1866_0,
c6288_wire_1866_1,
c6288_wire_1859_0,
c6288_wire_1859_1,
c6288_wire_1859_2,
c6288_wire_1862_0,
c6288_wire_1862_1,
c6288_wire_1870_0,
c6288_wire_1870_1,
c6288_wire_1875_0,
c6288_wire_1875_1,
c6288_wire_1880_0,
c6288_wire_1880_1,
c6288_wire_1885_0,
c6288_wire_1885_1,
c6288_wire_1891_0,
c6288_wire_1891_1,
c6288_wire_1897_0,
c6288_wire_1897_1,
c6288_wire_1902_0,
c6288_wire_1902_1,
c6288_wire_1907_0,
c6288_wire_1907_1,
c6288_wire_1912_0,
c6288_wire_1912_1,
c6288_wire_1917_0,
c6288_wire_1917_1,
c6288_wire_1922_0,
c6288_wire_1922_1,
c6288_wire_1927_0,
c6288_wire_1927_1,
c6288_wire_1867_0,
c6288_wire_1867_1,
c6288_wire_837_0,
c6288_wire_837_1,
c6288_wire_837_2,
c6288_wire_840_0,
c6288_wire_840_1,
c6288_wire_848_0,
c6288_wire_848_1,
c6288_wire_853_0,
c6288_wire_853_1,
c6288_wire_858_0,
c6288_wire_858_1,
c6288_wire_864_0,
c6288_wire_864_1,
c6288_wire_875_0,
c6288_wire_875_1,
c6288_wire_881_0,
c6288_wire_881_1,
c6288_wire_886_0,
c6288_wire_886_1,
c6288_wire_891_0,
c6288_wire_891_1,
c6288_wire_896_0,
c6288_wire_896_1,
c6288_wire_901_0,
c6288_wire_901_1,
c6288_wire_906_0,
c6288_wire_906_1,
c6288_wire_911_0,
c6288_wire_911_1,
c6288_wire_845_0,
c6288_wire_845_1,
c6288_wire_918_0,
c6288_wire_918_1,
c6288_wire_918_2,
c6288_wire_921_0,
c6288_wire_921_1,
c6288_wire_929_0,
c6288_wire_929_1,
c6288_wire_934_0,
c6288_wire_934_1,
c6288_wire_939_0,
c6288_wire_939_1,
c6288_wire_944_0,
c6288_wire_944_1,
c6288_wire_953_0,
c6288_wire_953_1,
c6288_wire_959_0,
c6288_wire_959_1,
c6288_wire_964_0,
c6288_wire_964_1,
c6288_wire_969_0,
c6288_wire_969_1,
c6288_wire_974_0,
c6288_wire_974_1,
c6288_wire_979_0,
c6288_wire_979_1,
c6288_wire_984_0,
c6288_wire_984_1,
c6288_wire_989_0,
c6288_wire_989_1,
c6288_wire_926_0,
c6288_wire_926_1,
c6288_wire_996_0,
c6288_wire_996_1,
c6288_wire_996_2,
c6288_wire_999_0,
c6288_wire_999_1,
c6288_wire_1007_0,
c6288_wire_1007_1,
c6288_wire_1012_0,
c6288_wire_1012_1,
c6288_wire_1017_0,
c6288_wire_1017_1,
c6288_wire_1022_0,
c6288_wire_1022_1,
c6288_wire_1031_0,
c6288_wire_1031_1,
c6288_wire_1037_0,
c6288_wire_1037_1,
c6288_wire_1042_0,
c6288_wire_1042_1,
c6288_wire_1047_0,
c6288_wire_1047_1,
c6288_wire_1052_0,
c6288_wire_1052_1,
c6288_wire_1057_0,
c6288_wire_1057_1,
c6288_wire_1062_0,
c6288_wire_1062_1,
c6288_wire_1067_0,
c6288_wire_1067_1,
c6288_wire_1004_0,
c6288_wire_1004_1,
c6288_wire_1073_0,
c6288_wire_1073_1,
c6288_wire_1075_0,
c6288_wire_1075_1,
c6288_wire_1083_0,
c6288_wire_1083_1,
c6288_wire_1088_0,
c6288_wire_1088_1,
c6288_wire_1093_0,
c6288_wire_1093_1,
c6288_wire_1098_0,
c6288_wire_1098_1,
c6288_wire_1109_0,
c6288_wire_1109_1,
c6288_wire_1109_2,
c6288_wire_1116_0,
c6288_wire_1116_1,
c6288_wire_1121_0,
c6288_wire_1121_1,
c6288_wire_1126_0,
c6288_wire_1126_1,
c6288_wire_1131_0,
c6288_wire_1131_1,
c6288_wire_1136_0,
c6288_wire_1136_1,
c6288_wire_1141_0,
c6288_wire_1141_1,
c6288_wire_1146_0,
c6288_wire_1146_1,
c6288_wire_1080_0,
c6288_wire_1080_1,
c6288_wire_746_0,
c6288_wire_746_1,
c6288_wire_746_2,
c6288_wire_750_0,
c6288_wire_750_1,
c6288_wire_759_0,
c6288_wire_759_1,
c6288_wire_765_0,
c6288_wire_765_1,
c6288_wire_771_0,
c6288_wire_771_1,
c6288_wire_777_0,
c6288_wire_777_1,
c6288_wire_786_0,
c6288_wire_786_1,
c6288_wire_793_0,
c6288_wire_793_1,
c6288_wire_799_0,
c6288_wire_799_1,
c6288_wire_805_0,
c6288_wire_805_1,
c6288_wire_811_0,
c6288_wire_811_1,
c6288_wire_817_0,
c6288_wire_817_1,
c6288_wire_823_0,
c6288_wire_823_1,
c6288_wire_829_0,
c6288_wire_829_1,
c6288_wire_755_0,
c6288_wire_755_1,
c6288_wire_1234_0,
c6288_wire_1234_1,
c6288_wire_1234_2,
c6288_wire_1237_0,
c6288_wire_1237_1,
c6288_wire_1245_0,
c6288_wire_1245_1,
c6288_wire_1250_0,
c6288_wire_1250_1,
c6288_wire_1255_0,
c6288_wire_1255_1,
c6288_wire_1260_0,
c6288_wire_1260_1,
c6288_wire_1270_0,
c6288_wire_1270_1,
c6288_wire_1276_0,
c6288_wire_1276_1,
c6288_wire_1281_0,
c6288_wire_1281_1,
c6288_wire_1286_0,
c6288_wire_1286_1,
c6288_wire_1291_0,
c6288_wire_1291_1,
c6288_wire_1296_0,
c6288_wire_1296_1,
c6288_wire_1301_0,
c6288_wire_1301_1,
c6288_wire_1306_0,
c6288_wire_1306_1,
c6288_wire_1242_0,
c6288_wire_1242_1,
c6288_wire_1313_0,
c6288_wire_1313_1,
c6288_wire_1313_2,
c6288_wire_1316_0,
c6288_wire_1316_1,
c6288_wire_1324_0,
c6288_wire_1324_1,
c6288_wire_1329_0,
c6288_wire_1329_1,
c6288_wire_1334_0,
c6288_wire_1334_1,
c6288_wire_1339_0,
c6288_wire_1339_1,
c6288_wire_1348_0,
c6288_wire_1348_1,
c6288_wire_1354_0,
c6288_wire_1354_1,
c6288_wire_1359_0,
c6288_wire_1359_1,
c6288_wire_1364_0,
c6288_wire_1364_1,
c6288_wire_1369_0,
c6288_wire_1369_1,
c6288_wire_1374_0,
c6288_wire_1374_1,
c6288_wire_1379_0,
c6288_wire_1379_1,
c6288_wire_1384_0,
c6288_wire_1384_1,
c6288_wire_1321_0,
c6288_wire_1321_1,
c6288_wire_1391_0,
c6288_wire_1391_1,
c6288_wire_1391_2,
c6288_wire_1394_0,
c6288_wire_1394_1,
c6288_wire_1402_0,
c6288_wire_1402_1,
c6288_wire_1407_0,
c6288_wire_1407_1,
c6288_wire_1412_0,
c6288_wire_1412_1,
c6288_wire_1417_0,
c6288_wire_1417_1,
c6288_wire_1426_0,
c6288_wire_1426_1,
c6288_wire_1432_0,
c6288_wire_1432_1,
c6288_wire_1437_0,
c6288_wire_1437_1,
c6288_wire_1442_0,
c6288_wire_1442_1,
c6288_wire_1447_0,
c6288_wire_1447_1,
c6288_wire_1452_0,
c6288_wire_1452_1,
c6288_wire_1457_0,
c6288_wire_1457_1,
c6288_wire_1462_0,
c6288_wire_1462_1,
c6288_wire_1399_0,
c6288_wire_1399_1,
c6288_wire_1469_0,
c6288_wire_1469_1,
c6288_wire_1469_2,
c6288_wire_1472_0,
c6288_wire_1472_1,
c6288_wire_1480_0,
c6288_wire_1480_1,
c6288_wire_1485_0,
c6288_wire_1485_1,
c6288_wire_1490_0,
c6288_wire_1490_1,
c6288_wire_1495_0,
c6288_wire_1495_1,
c6288_wire_1504_0,
c6288_wire_1504_1,
c6288_wire_1510_0,
c6288_wire_1510_1,
c6288_wire_1515_0,
c6288_wire_1515_1,
c6288_wire_1520_0,
c6288_wire_1520_1,
c6288_wire_1525_0,
c6288_wire_1525_1,
c6288_wire_1530_0,
c6288_wire_1530_1,
c6288_wire_1535_0,
c6288_wire_1535_1,
c6288_wire_1540_0,
c6288_wire_1540_1,
c6288_wire_1477_0,
c6288_wire_1477_1,
c6288_wire_1547_0,
c6288_wire_1547_1,
c6288_wire_1547_2,
c6288_wire_1550_0,
c6288_wire_1550_1,
c6288_wire_1558_0,
c6288_wire_1558_1,
c6288_wire_1563_0,
c6288_wire_1563_1,
c6288_wire_1568_0,
c6288_wire_1568_1,
c6288_wire_1573_0,
c6288_wire_1573_1,
c6288_wire_1582_0,
c6288_wire_1582_1,
c6288_wire_1588_0,
c6288_wire_1588_1,
c6288_wire_1593_0,
c6288_wire_1593_1,
c6288_wire_1598_0,
c6288_wire_1598_1,
c6288_wire_1603_0,
c6288_wire_1603_1,
c6288_wire_1608_0,
c6288_wire_1608_1,
c6288_wire_1613_0,
c6288_wire_1613_1,
c6288_wire_1618_0,
c6288_wire_1618_1,
c6288_wire_1555_0,
c6288_wire_1555_1,
c6288_wire_1625_0,
c6288_wire_1625_1,
c6288_wire_1625_2,
c6288_wire_1628_0,
c6288_wire_1628_1,
c6288_wire_1636_0,
c6288_wire_1636_1,
c6288_wire_1641_0,
c6288_wire_1641_1,
c6288_wire_1646_0,
c6288_wire_1646_1,
c6288_wire_1651_0,
c6288_wire_1651_1,
c6288_wire_1660_0,
c6288_wire_1660_1,
c6288_wire_1666_0,
c6288_wire_1666_1,
c6288_wire_1671_0,
c6288_wire_1671_1,
c6288_wire_1676_0,
c6288_wire_1676_1,
c6288_wire_1681_0,
c6288_wire_1681_1,
c6288_wire_1686_0,
c6288_wire_1686_1,
c6288_wire_1691_0,
c6288_wire_1691_1,
c6288_wire_1696_0,
c6288_wire_1696_1,
c6288_wire_1633_0,
c6288_wire_1633_1,
c6288_wire_1703_0,
c6288_wire_1703_1,
c6288_wire_1703_2,
c6288_wire_1706_0,
c6288_wire_1706_1,
c6288_wire_1714_0,
c6288_wire_1714_1,
c6288_wire_1719_0,
c6288_wire_1719_1,
c6288_wire_1724_0,
c6288_wire_1724_1,
c6288_wire_1729_0,
c6288_wire_1729_1,
c6288_wire_1738_0,
c6288_wire_1738_1,
c6288_wire_1744_0,
c6288_wire_1744_1,
c6288_wire_1749_0,
c6288_wire_1749_1,
c6288_wire_1754_0,
c6288_wire_1754_1,
c6288_wire_1759_0,
c6288_wire_1759_1,
c6288_wire_1764_0,
c6288_wire_1764_1,
c6288_wire_1769_0,
c6288_wire_1769_1,
c6288_wire_1774_0,
c6288_wire_1774_1,
c6288_wire_1711_0,
c6288_wire_1711_1,
c6288_wire_1781_0,
c6288_wire_1781_1,
c6288_wire_1781_2,
c6288_wire_1784_0,
c6288_wire_1784_1,
c6288_wire_1792_0,
c6288_wire_1792_1,
c6288_wire_1797_0,
c6288_wire_1797_1,
c6288_wire_1802_0,
c6288_wire_1802_1,
c6288_wire_1807_0,
c6288_wire_1807_1,
c6288_wire_1816_0,
c6288_wire_1816_1,
c6288_wire_1822_0,
c6288_wire_1822_1,
c6288_wire_1827_0,
c6288_wire_1827_1,
c6288_wire_1832_0,
c6288_wire_1832_1,
c6288_wire_1837_0,
c6288_wire_1837_1,
c6288_wire_1842_0,
c6288_wire_1842_1,
c6288_wire_1847_0,
c6288_wire_1847_1,
c6288_wire_1852_0,
c6288_wire_1852_1,
c6288_wire_1789_0,
c6288_wire_1789_1,
c6288_wire_2015_0,
c6288_wire_2015_1,
c6288_wire_2015_2,
c6288_wire_160_0,
c6288_wire_160_1,
c6288_wire_160_2,
c6288_wire_202_0,
c6288_wire_202_1,
c6288_wire_202_2,
c6288_wire_244_0,
c6288_wire_244_1,
c6288_wire_244_2,
c6288_wire_284_0,
c6288_wire_284_1,
c6288_wire_284_2,
c6288_wire_311_0,
c6288_wire_311_1,
c6288_wire_311_2,
c6288_wire_309_0,
c6288_wire_309_1,
c6288_wire_309_2,
c6288_wire_307_0,
c6288_wire_307_1,
c6288_wire_307_2,
c6288_wire_305_0,
c6288_wire_305_1,
c6288_wire_305_2,
c6288_wire_303_0,
c6288_wire_303_1,
c6288_wire_303_2,
c6288_wire_1104_0,
c6288_wire_1104_1,
c6288_wire_2230_0,
c6288_wire_2230_1,
c6288_wire_2230_2,
c6288_wire_325_0,
c6288_wire_325_1,
c6288_wire_325_2,
c6288_wire_323_0,
c6288_wire_323_1,
c6288_wire_323_2,
c6288_wire_321_0,
c6288_wire_321_1,
c6288_wire_321_2,
c6288_wire_319_0,
c6288_wire_319_1,
c6288_wire_319_2,
c6288_wire_317_0,
c6288_wire_317_1,
c6288_wire_317_2,
c6288_wire_315_0,
c6288_wire_315_1,
c6288_wire_315_2,
c6288_wire_313_0,
c6288_wire_313_1,
c6288_wire_313_2,
c6288_wire_402_0,
c6288_wire_402_1,
c6288_wire_402_2,
c6288_wire_444_0,
c6288_wire_444_1,
c6288_wire_444_2,
c6288_wire_486_0,
c6288_wire_486_1,
c6288_wire_486_2,
c6288_wire_528_0,
c6288_wire_528_1,
c6288_wire_528_2,
c6288_wire_570_0,
c6288_wire_570_1,
c6288_wire_570_2,
c6288_wire_612_0,
c6288_wire_612_1,
c6288_wire_612_2,
c6288_wire_654_0,
c6288_wire_654_1,
c6288_wire_654_2,
c6288_wire_696_0,
c6288_wire_696_1,
c6288_wire_696_2,
c6288_wire_738_0,
c6288_wire_738_1,
c6288_wire_738_2,
c6288_wire_756_0,
c6288_wire_756_1,
c6288_wire_762_0,
c6288_wire_762_1,
c6288_wire_768_0,
c6288_wire_768_1,
c6288_wire_774_0,
c6288_wire_774_1,
c6288_wire_779_0,
c6288_wire_779_1,
c6288_wire_790_0,
c6288_wire_790_1,
c6288_wire_796_0,
c6288_wire_796_1,
c6288_wire_802_0,
c6288_wire_802_1,
c6288_wire_808_0,
c6288_wire_808_1,
c6288_wire_814_0,
c6288_wire_814_1,
c6288_wire_820_0,
c6288_wire_820_1,
c6288_wire_826_0,
c6288_wire_826_1,
c6288_wire_832_0,
c6288_wire_832_1,
c6288_wire_835_0,
c6288_wire_835_1,
c6288_wire_740_0,
c6288_wire_740_1,
c6288_wire_740_2,
c6288_wire_740_3,
c6288_wire_32_0,
c6288_wire_32_1,
c6288_wire_32_2,
c6288_wire_32_3,
c6288_wire_32_4,
c6288_wire_32_5,
c6288_wire_32_6,
c6288_wire_32_7,
c6288_wire_32_8,
c6288_wire_32_9,
c6288_wire_32_10,
c6288_wire_32_11,
c6288_wire_32_12,
c6288_wire_32_13,
c6288_wire_32_14,
c6288_wire_32_15,
c6288_wire_32_16,
c6288_wire_32_17,
c6288_wire_32_18,
c6288_wire_32_19,
c6288_wire_32_20,
c6288_wire_32_21,
c6288_wire_32_22,
c6288_wire_32_23,
c6288_wire_32_24,
c6288_wire_32_25,
c6288_wire_32_26,
c6288_wire_32_27,
c6288_wire_32_28,
c6288_wire_32_29,
c6288_wire_32_30,
c6288_wire_32_31,
c6288_wire_57_0,
c6288_wire_57_1,
c6288_wire_57_2,
c6288_wire_57_3,
c6288_wire_57_4,
c6288_wire_57_5,
c6288_wire_57_6,
c6288_wire_57_7,
c6288_wire_57_8,
c6288_wire_57_9,
c6288_wire_57_10,
c6288_wire_57_11,
c6288_wire_57_12,
c6288_wire_57_13,
c6288_wire_57_14,
c6288_wire_57_15,
c6288_wire_57_16,
c6288_wire_57_17,
c6288_wire_57_18,
c6288_wire_57_19,
c6288_wire_57_20,
c6288_wire_57_21,
c6288_wire_57_22,
c6288_wire_57_23,
c6288_wire_57_24,
c6288_wire_57_25,
c6288_wire_57_26,
c6288_wire_57_27,
c6288_wire_57_28,
c6288_wire_57_29,
c6288_wire_57_30,
c6288_wire_57_31,
c6288_wire_57_32,
c6288_wire_57_33,
c6288_wire_57_34,
c6288_wire_57_35,
c6288_wire_57_36,
c6288_wire_57_37,
c6288_wire_57_38,
c6288_wire_57_39,
c6288_wire_57_40,
c6288_wire_57_41,
c6288_wire_57_42,
c6288_wire_57_43,
c6288_wire_57_44,
c6288_wire_57_45,
c6288_wire_62_0,
c6288_wire_62_1,
c6288_wire_62_2,
c6288_wire_62_3,
c6288_wire_62_4,
c6288_wire_62_5,
c6288_wire_62_6,
c6288_wire_62_7,
c6288_wire_62_8,
c6288_wire_62_9,
c6288_wire_62_10,
c6288_wire_62_11,
c6288_wire_62_12,
c6288_wire_62_13,
c6288_wire_62_14,
c6288_wire_62_15,
c6288_wire_62_16,
c6288_wire_62_17,
c6288_wire_62_18,
c6288_wire_62_19,
c6288_wire_62_20,
c6288_wire_62_21,
c6288_wire_62_22,
c6288_wire_62_23,
c6288_wire_62_24,
c6288_wire_62_25,
c6288_wire_62_26,
c6288_wire_62_27,
c6288_wire_62_28,
c6288_wire_62_29,
c6288_wire_62_30,
c6288_wire_62_31,
c6288_wire_62_32,
c6288_wire_62_33,
c6288_wire_62_34,
c6288_wire_62_35,
c6288_wire_62_36,
c6288_wire_62_37,
c6288_wire_62_38,
c6288_wire_62_39,
c6288_wire_62_40,
c6288_wire_62_41,
c6288_wire_62_42,
c6288_wire_62_43,
c6288_wire_62_44,
c6288_wire_62_45,
c6288_wire_67_0,
c6288_wire_67_1,
c6288_wire_67_2,
c6288_wire_67_3,
c6288_wire_67_4,
c6288_wire_67_5,
c6288_wire_67_6,
c6288_wire_67_7,
c6288_wire_67_8,
c6288_wire_67_9,
c6288_wire_67_10,
c6288_wire_67_11,
c6288_wire_67_12,
c6288_wire_67_13,
c6288_wire_67_14,
c6288_wire_67_15,
c6288_wire_67_16,
c6288_wire_67_17,
c6288_wire_67_18,
c6288_wire_67_19,
c6288_wire_67_20,
c6288_wire_67_21,
c6288_wire_67_22,
c6288_wire_67_23,
c6288_wire_67_24,
c6288_wire_67_25,
c6288_wire_67_26,
c6288_wire_67_27,
c6288_wire_67_28,
c6288_wire_67_29,
c6288_wire_67_30,
c6288_wire_67_31,
c6288_wire_67_32,
c6288_wire_67_33,
c6288_wire_67_34,
c6288_wire_67_35,
c6288_wire_67_36,
c6288_wire_67_37,
c6288_wire_67_38,
c6288_wire_67_39,
c6288_wire_67_40,
c6288_wire_67_41,
c6288_wire_67_42,
c6288_wire_67_43,
c6288_wire_67_44,
c6288_wire_67_45,
c6288_wire_5_0,
c6288_wire_5_1,
c6288_wire_5_2,
c6288_wire_5_3,
c6288_wire_5_4,
c6288_wire_5_5,
c6288_wire_5_6,
c6288_wire_5_7,
c6288_wire_5_8,
c6288_wire_5_9,
c6288_wire_5_10,
c6288_wire_5_11,
c6288_wire_5_12,
c6288_wire_5_13,
c6288_wire_5_14,
c6288_wire_5_15,
c6288_wire_5_16,
c6288_wire_5_17,
c6288_wire_5_18,
c6288_wire_5_19,
c6288_wire_5_20,
c6288_wire_5_21,
c6288_wire_5_22,
c6288_wire_5_23,
c6288_wire_5_24,
c6288_wire_5_25,
c6288_wire_5_26,
c6288_wire_5_27,
c6288_wire_5_28,
c6288_wire_5_29,
c6288_wire_5_30,
c6288_wire_5_31,
c6288_wire_5_32,
c6288_wire_5_33,
c6288_wire_5_34,
c6288_wire_5_35,
c6288_wire_5_36,
c6288_wire_5_37,
c6288_wire_5_38,
c6288_wire_5_39,
c6288_wire_5_40,
c6288_wire_5_41,
c6288_wire_5_42,
c6288_wire_5_43,
c6288_wire_5_44,
c6288_wire_5_45,
c6288_wire_2_0,
c6288_wire_2_1,
c6288_wire_2_2,
c6288_wire_2_3,
c6288_wire_2_4,
c6288_wire_2_5,
c6288_wire_2_6,
c6288_wire_2_7,
c6288_wire_2_8,
c6288_wire_2_9,
c6288_wire_2_10,
c6288_wire_2_11,
c6288_wire_2_12,
c6288_wire_2_13,
c6288_wire_2_14,
c6288_wire_2_15,
c6288_wire_2_16,
c6288_wire_2_17,
c6288_wire_2_18,
c6288_wire_2_19,
c6288_wire_2_20,
c6288_wire_2_21,
c6288_wire_2_22,
c6288_wire_2_23,
c6288_wire_2_24,
c6288_wire_2_25,
c6288_wire_2_26,
c6288_wire_2_27,
c6288_wire_2_28,
c6288_wire_2_29,
c6288_wire_2_30,
c6288_wire_2_31,
c6288_wire_2_32,
c6288_wire_2_33,
c6288_wire_2_34,
c6288_wire_2_35,
c6288_wire_2_36,
c6288_wire_2_37,
c6288_wire_2_38,
c6288_wire_2_39,
c6288_wire_2_40,
c6288_wire_2_41,
c6288_wire_2_42,
c6288_wire_2_43,
c6288_wire_2_44,
c6288_wire_2_45,
c6288_wire_30_0,
c6288_wire_30_1,
c6288_wire_30_2,
c6288_wire_30_3,
c6288_wire_30_4,
c6288_wire_30_5,
c6288_wire_30_6,
c6288_wire_30_7,
c6288_wire_30_8,
c6288_wire_30_9,
c6288_wire_30_10,
c6288_wire_30_11,
c6288_wire_30_12,
c6288_wire_30_13,
c6288_wire_30_14,
c6288_wire_30_15,
c6288_wire_30_16,
c6288_wire_30_17,
c6288_wire_30_18,
c6288_wire_30_19,
c6288_wire_30_20,
c6288_wire_30_21,
c6288_wire_30_22,
c6288_wire_30_23,
c6288_wire_30_24,
c6288_wire_30_25,
c6288_wire_30_26,
c6288_wire_30_27,
c6288_wire_30_28,
c6288_wire_30_29,
c6288_wire_30_30,
c6288_wire_30_31,
c6288_wire_30_32,
c6288_wire_30_33,
c6288_wire_30_34,
c6288_wire_30_35,
c6288_wire_30_36,
c6288_wire_30_37,
c6288_wire_30_38,
c6288_wire_30_39,
c6288_wire_30_40,
c6288_wire_30_41,
c6288_wire_30_42,
c6288_wire_30_43,
c6288_wire_30_44,
c6288_wire_30_45,
c6288_wire_10_0,
c6288_wire_10_1,
c6288_wire_10_2,
c6288_wire_10_3,
c6288_wire_10_4,
c6288_wire_10_5,
c6288_wire_10_6,
c6288_wire_10_7,
c6288_wire_10_8,
c6288_wire_10_9,
c6288_wire_10_10,
c6288_wire_10_11,
c6288_wire_10_12,
c6288_wire_10_13,
c6288_wire_10_14,
c6288_wire_10_15,
c6288_wire_10_16,
c6288_wire_10_17,
c6288_wire_10_18,
c6288_wire_10_19,
c6288_wire_10_20,
c6288_wire_10_21,
c6288_wire_10_22,
c6288_wire_10_23,
c6288_wire_10_24,
c6288_wire_10_25,
c6288_wire_10_26,
c6288_wire_10_27,
c6288_wire_10_28,
c6288_wire_10_29,
c6288_wire_10_30,
c6288_wire_10_31,
c6288_wire_10_32,
c6288_wire_10_33,
c6288_wire_10_34,
c6288_wire_10_35,
c6288_wire_10_36,
c6288_wire_10_37,
c6288_wire_10_38,
c6288_wire_10_39,
c6288_wire_10_40,
c6288_wire_10_41,
c6288_wire_10_42,
c6288_wire_10_43,
c6288_wire_10_44,
c6288_wire_10_45,
c6288_wire_15_0,
c6288_wire_15_1,
c6288_wire_15_2,
c6288_wire_15_3,
c6288_wire_15_4,
c6288_wire_15_5,
c6288_wire_15_6,
c6288_wire_15_7,
c6288_wire_15_8,
c6288_wire_15_9,
c6288_wire_15_10,
c6288_wire_15_11,
c6288_wire_15_12,
c6288_wire_15_13,
c6288_wire_15_14,
c6288_wire_15_15,
c6288_wire_15_16,
c6288_wire_15_17,
c6288_wire_15_18,
c6288_wire_15_19,
c6288_wire_15_20,
c6288_wire_15_21,
c6288_wire_15_22,
c6288_wire_15_23,
c6288_wire_15_24,
c6288_wire_15_25,
c6288_wire_15_26,
c6288_wire_15_27,
c6288_wire_15_28,
c6288_wire_15_29,
c6288_wire_15_30,
c6288_wire_15_31,
c6288_wire_15_32,
c6288_wire_15_33,
c6288_wire_15_34,
c6288_wire_15_35,
c6288_wire_15_36,
c6288_wire_15_37,
c6288_wire_15_38,
c6288_wire_15_39,
c6288_wire_15_40,
c6288_wire_15_41,
c6288_wire_15_42,
c6288_wire_15_43,
c6288_wire_15_44,
c6288_wire_15_45,
c6288_wire_20_0,
c6288_wire_20_1,
c6288_wire_20_2,
c6288_wire_20_3,
c6288_wire_20_4,
c6288_wire_20_5,
c6288_wire_20_6,
c6288_wire_20_7,
c6288_wire_20_8,
c6288_wire_20_9,
c6288_wire_20_10,
c6288_wire_20_11,
c6288_wire_20_12,
c6288_wire_20_13,
c6288_wire_20_14,
c6288_wire_20_15,
c6288_wire_20_16,
c6288_wire_20_17,
c6288_wire_20_18,
c6288_wire_20_19,
c6288_wire_20_20,
c6288_wire_20_21,
c6288_wire_20_22,
c6288_wire_20_23,
c6288_wire_20_24,
c6288_wire_20_25,
c6288_wire_20_26,
c6288_wire_20_27,
c6288_wire_20_28,
c6288_wire_20_29,
c6288_wire_20_30,
c6288_wire_20_31,
c6288_wire_20_32,
c6288_wire_20_33,
c6288_wire_20_34,
c6288_wire_20_35,
c6288_wire_20_36,
c6288_wire_20_37,
c6288_wire_20_38,
c6288_wire_20_39,
c6288_wire_20_40,
c6288_wire_20_41,
c6288_wire_20_42,
c6288_wire_20_43,
c6288_wire_20_44,
c6288_wire_20_45,
c6288_wire_25_0,
c6288_wire_25_1,
c6288_wire_25_2,
c6288_wire_25_3,
c6288_wire_25_4,
c6288_wire_25_5,
c6288_wire_25_6,
c6288_wire_25_7,
c6288_wire_25_8,
c6288_wire_25_9,
c6288_wire_25_10,
c6288_wire_25_11,
c6288_wire_25_12,
c6288_wire_25_13,
c6288_wire_25_14,
c6288_wire_25_15,
c6288_wire_25_16,
c6288_wire_25_17,
c6288_wire_25_18,
c6288_wire_25_19,
c6288_wire_25_20,
c6288_wire_25_21,
c6288_wire_25_22,
c6288_wire_25_23,
c6288_wire_25_24,
c6288_wire_25_25,
c6288_wire_25_26,
c6288_wire_25_27,
c6288_wire_25_28,
c6288_wire_25_29,
c6288_wire_25_30,
c6288_wire_25_31,
c6288_wire_25_32,
c6288_wire_25_33,
c6288_wire_25_34,
c6288_wire_25_35,
c6288_wire_25_36,
c6288_wire_25_37,
c6288_wire_25_38,
c6288_wire_25_39,
c6288_wire_25_40,
c6288_wire_25_41,
c6288_wire_25_42,
c6288_wire_25_43,
c6288_wire_25_44,
c6288_wire_330_0,
c6288_wire_330_1,
c6288_wire_330_2,
c6288_wire_330_3,
c6288_wire_330_4,
c6288_wire_330_5,
c6288_wire_330_6,
c6288_wire_330_7,
c6288_wire_330_8,
c6288_wire_330_9,
c6288_wire_330_10,
c6288_wire_330_11,
c6288_wire_330_12,
c6288_wire_330_13,
c6288_wire_330_14,
c6288_wire_330_15,
c6288_wire_330_16,
c6288_wire_330_17,
c6288_wire_330_18,
c6288_wire_330_19,
c6288_wire_330_20,
c6288_wire_330_21,
c6288_wire_330_22,
c6288_wire_330_23,
c6288_wire_330_24,
c6288_wire_330_25,
c6288_wire_330_26,
c6288_wire_330_27,
c6288_wire_330_28,
c6288_wire_330_29,
c6288_wire_330_30,
c6288_wire_330_31,
c6288_wire_330_32,
c6288_wire_330_33,
c6288_wire_330_34,
c6288_wire_330_35,
c6288_wire_330_36,
c6288_wire_330_37,
c6288_wire_330_38,
c6288_wire_330_39,
c6288_wire_330_40,
c6288_wire_330_41,
c6288_wire_330_42,
c6288_wire_330_43,
c6288_wire_3_0,
c6288_wire_3_1,
c6288_wire_3_2,
c6288_wire_3_3,
c6288_wire_3_4,
c6288_wire_3_5,
c6288_wire_3_6,
c6288_wire_3_7,
c6288_wire_3_8,
c6288_wire_3_9,
c6288_wire_3_10,
c6288_wire_3_11,
c6288_wire_3_12,
c6288_wire_3_13,
c6288_wire_3_14,
c6288_wire_3_15,
c6288_wire_3_16,
c6288_wire_3_17,
c6288_wire_6_0,
c6288_wire_6_1,
c6288_wire_6_2,
c6288_wire_6_3,
c6288_wire_6_4,
c6288_wire_6_5,
c6288_wire_6_6,
c6288_wire_6_7,
c6288_wire_6_8,
c6288_wire_6_9,
c6288_wire_6_10,
c6288_wire_6_11,
c6288_wire_6_12,
c6288_wire_6_13,
c6288_wire_6_14,
c6288_wire_6_15,
c6288_wire_6_16,
c6288_wire_6_17,
c6288_wire_6_18,
c6288_wire_6_19,
c6288_wire_6_20,
c6288_wire_6_21,
c6288_wire_6_22,
c6288_wire_6_23,
c6288_wire_6_24,
c6288_wire_6_25,
c6288_wire_6_26,
c6288_wire_6_27,
c6288_wire_6_28,
c6288_wire_6_29,
c6288_wire_6_30,
c6288_wire_6_31,
c6288_wire_6_32,
c6288_wire_6_33,
c6288_wire_6_34,
c6288_wire_6_35,
c6288_wire_6_36,
c6288_wire_6_37,
c6288_wire_6_38,
c6288_wire_6_39,
c6288_wire_6_40,
c6288_wire_6_41,
c6288_wire_6_42,
c6288_wire_6_43,
c6288_wire_6_44,
c6288_wire_6_45,
c6288_wire_6_46,
c6288_wire_6_47,
c6288_wire_78_0,
c6288_wire_78_1,
c6288_wire_78_2,
c6288_wire_78_3,
c6288_wire_78_4,
c6288_wire_78_5,
c6288_wire_78_6,
c6288_wire_78_7,
c6288_wire_78_8,
c6288_wire_78_9,
c6288_wire_78_10,
c6288_wire_78_11,
c6288_wire_78_12,
c6288_wire_78_13,
c6288_wire_78_14,
c6288_wire_78_15,
c6288_wire_78_16,
c6288_wire_78_17,
c6288_wire_78_18,
c6288_wire_78_19,
c6288_wire_78_20,
c6288_wire_78_21,
c6288_wire_78_22,
c6288_wire_78_23,
c6288_wire_78_24,
c6288_wire_78_25,
c6288_wire_78_26,
c6288_wire_78_27,
c6288_wire_78_28,
c6288_wire_78_29,
c6288_wire_78_30,
c6288_wire_78_31,
c6288_wire_78_32,
c6288_wire_78_33,
c6288_wire_78_34,
c6288_wire_78_35,
c6288_wire_78_36,
c6288_wire_78_37,
c6288_wire_78_38,
c6288_wire_78_39,
c6288_wire_78_40,
c6288_wire_78_41,
c6288_wire_78_42,
c6288_wire_78_43,
c6288_wire_78_44,
c6288_wire_78_45,
c6288_wire_81_0,
c6288_wire_81_1,
c6288_wire_81_2,
c6288_wire_81_3,
c6288_wire_81_4,
c6288_wire_81_5,
c6288_wire_81_6,
c6288_wire_81_7,
c6288_wire_81_8,
c6288_wire_81_9,
c6288_wire_81_10,
c6288_wire_81_11,
c6288_wire_81_12,
c6288_wire_81_13,
c6288_wire_81_14,
c6288_wire_81_15,
c6288_wire_81_16,
c6288_wire_81_17,
c6288_wire_81_18,
c6288_wire_81_19,
c6288_wire_81_20,
c6288_wire_81_21,
c6288_wire_81_22,
c6288_wire_81_23,
c6288_wire_81_24,
c6288_wire_81_25,
c6288_wire_81_26,
c6288_wire_81_27,
c6288_wire_81_28,
c6288_wire_81_29,
c6288_wire_81_30,
c6288_wire_81_31,
c6288_wire_81_32,
c6288_wire_81_33,
c6288_wire_81_34,
c6288_wire_81_35,
c6288_wire_81_36,
c6288_wire_81_37,
c6288_wire_81_38,
c6288_wire_81_39,
c6288_wire_81_40,
c6288_wire_81_41,
c6288_wire_81_42,
c6288_wire_81_43,
c6288_wire_81_44,
c6288_wire_81_45,
c6288_wire_81_46,
c6288_wire_84_0,
c6288_wire_84_1,
c6288_wire_84_2,
c6288_wire_84_3,
c6288_wire_84_4,
c6288_wire_84_5,
c6288_wire_84_6,
c6288_wire_84_7,
c6288_wire_84_8,
c6288_wire_84_9,
c6288_wire_84_10,
c6288_wire_84_11,
c6288_wire_84_12,
c6288_wire_84_13,
c6288_wire_84_14,
c6288_wire_84_15,
c6288_wire_84_16,
c6288_wire_84_17,
c6288_wire_84_18,
c6288_wire_84_19,
c6288_wire_84_20,
c6288_wire_84_21,
c6288_wire_84_22,
c6288_wire_84_23,
c6288_wire_84_24,
c6288_wire_84_25,
c6288_wire_84_26,
c6288_wire_84_27,
c6288_wire_84_28,
c6288_wire_84_29,
c6288_wire_84_30,
c6288_wire_84_31,
c6288_wire_84_32,
c6288_wire_84_33,
c6288_wire_84_34,
c6288_wire_84_35,
c6288_wire_84_36,
c6288_wire_84_37,
c6288_wire_84_38,
c6288_wire_84_39,
c6288_wire_84_40,
c6288_wire_84_41,
c6288_wire_84_42,
c6288_wire_84_43,
c6288_wire_84_44,
c6288_wire_84_45,
c6288_wire_84_46,
c6288_wire_37_0,
c6288_wire_37_1,
c6288_wire_37_2,
c6288_wire_37_3,
c6288_wire_37_4,
c6288_wire_37_5,
c6288_wire_37_6,
c6288_wire_37_7,
c6288_wire_37_8,
c6288_wire_37_9,
c6288_wire_37_10,
c6288_wire_37_11,
c6288_wire_37_12,
c6288_wire_37_13,
c6288_wire_37_14,
c6288_wire_37_15,
c6288_wire_37_16,
c6288_wire_37_17,
c6288_wire_37_18,
c6288_wire_37_19,
c6288_wire_37_20,
c6288_wire_37_21,
c6288_wire_37_22,
c6288_wire_37_23,
c6288_wire_37_24,
c6288_wire_37_25,
c6288_wire_37_26,
c6288_wire_37_27,
c6288_wire_37_28,
c6288_wire_37_29,
c6288_wire_37_30,
c6288_wire_37_31,
c6288_wire_37_32,
c6288_wire_37_33,
c6288_wire_37_34,
c6288_wire_37_35,
c6288_wire_37_36,
c6288_wire_37_37,
c6288_wire_37_38,
c6288_wire_37_39,
c6288_wire_37_40,
c6288_wire_37_41,
c6288_wire_37_42,
c6288_wire_37_43,
c6288_wire_37_44,
c6288_wire_37_45,
c6288_wire_87_0,
c6288_wire_87_1,
c6288_wire_87_2,
c6288_wire_87_3,
c6288_wire_87_4,
c6288_wire_87_5,
c6288_wire_87_6,
c6288_wire_87_7,
c6288_wire_87_8,
c6288_wire_87_9,
c6288_wire_87_10,
c6288_wire_87_11,
c6288_wire_87_12,
c6288_wire_87_13,
c6288_wire_87_14,
c6288_wire_87_15,
c6288_wire_87_16,
c6288_wire_87_17,
c6288_wire_87_18,
c6288_wire_87_19,
c6288_wire_87_20,
c6288_wire_87_21,
c6288_wire_87_22,
c6288_wire_87_23,
c6288_wire_87_24,
c6288_wire_87_25,
c6288_wire_87_26,
c6288_wire_87_27,
c6288_wire_87_28,
c6288_wire_87_29,
c6288_wire_87_30,
c6288_wire_87_31,
c6288_wire_87_32,
c6288_wire_87_33,
c6288_wire_87_34,
c6288_wire_87_35,
c6288_wire_87_36,
c6288_wire_87_37,
c6288_wire_87_38,
c6288_wire_87_39,
c6288_wire_87_40,
c6288_wire_87_41,
c6288_wire_87_42,
c6288_wire_87_43,
c6288_wire_87_44,
c6288_wire_87_45,
c6288_wire_87_46,
c6288_wire_90_0,
c6288_wire_90_1,
c6288_wire_90_2,
c6288_wire_90_3,
c6288_wire_90_4,
c6288_wire_90_5,
c6288_wire_90_6,
c6288_wire_90_7,
c6288_wire_90_8,
c6288_wire_90_9,
c6288_wire_90_10,
c6288_wire_90_11,
c6288_wire_90_12,
c6288_wire_90_13,
c6288_wire_90_14,
c6288_wire_90_15,
c6288_wire_90_16,
c6288_wire_90_17,
c6288_wire_90_18,
c6288_wire_90_19,
c6288_wire_90_20,
c6288_wire_90_21,
c6288_wire_90_22,
c6288_wire_90_23,
c6288_wire_90_24,
c6288_wire_90_25,
c6288_wire_90_26,
c6288_wire_90_27,
c6288_wire_90_28,
c6288_wire_90_29,
c6288_wire_90_30,
c6288_wire_90_31,
c6288_wire_90_32,
c6288_wire_90_33,
c6288_wire_90_34,
c6288_wire_90_35,
c6288_wire_90_36,
c6288_wire_90_37,
c6288_wire_90_38,
c6288_wire_90_39,
c6288_wire_90_40,
c6288_wire_90_41,
c6288_wire_90_42,
c6288_wire_90_43,
c6288_wire_90_44,
c6288_wire_90_45,
c6288_wire_90_46,
c6288_wire_93_0,
c6288_wire_93_1,
c6288_wire_93_2,
c6288_wire_93_3,
c6288_wire_93_4,
c6288_wire_93_5,
c6288_wire_93_6,
c6288_wire_93_7,
c6288_wire_93_8,
c6288_wire_93_9,
c6288_wire_93_10,
c6288_wire_93_11,
c6288_wire_93_12,
c6288_wire_93_13,
c6288_wire_93_14,
c6288_wire_93_15,
c6288_wire_93_16,
c6288_wire_93_17,
c6288_wire_93_18,
c6288_wire_93_19,
c6288_wire_93_20,
c6288_wire_93_21,
c6288_wire_93_22,
c6288_wire_93_23,
c6288_wire_93_24,
c6288_wire_93_25,
c6288_wire_93_26,
c6288_wire_93_27,
c6288_wire_93_28,
c6288_wire_93_29,
c6288_wire_93_30,
c6288_wire_93_31,
c6288_wire_93_32,
c6288_wire_93_33,
c6288_wire_93_34,
c6288_wire_93_35,
c6288_wire_93_36,
c6288_wire_93_37,
c6288_wire_93_38,
c6288_wire_93_39,
c6288_wire_93_40,
c6288_wire_93_41,
c6288_wire_93_42,
c6288_wire_93_43,
c6288_wire_93_44,
c6288_wire_93_45,
c6288_wire_93_46,
c6288_wire_96_0,
c6288_wire_96_1,
c6288_wire_96_2,
c6288_wire_96_3,
c6288_wire_96_4,
c6288_wire_96_5,
c6288_wire_96_6,
c6288_wire_96_7,
c6288_wire_96_8,
c6288_wire_96_9,
c6288_wire_96_10,
c6288_wire_96_11,
c6288_wire_96_12,
c6288_wire_96_13,
c6288_wire_96_14,
c6288_wire_96_15,
c6288_wire_96_16,
c6288_wire_96_17,
c6288_wire_96_18,
c6288_wire_96_19,
c6288_wire_96_20,
c6288_wire_96_21,
c6288_wire_96_22,
c6288_wire_96_23,
c6288_wire_96_24,
c6288_wire_96_25,
c6288_wire_96_26,
c6288_wire_96_27,
c6288_wire_96_28,
c6288_wire_96_29,
c6288_wire_96_30,
c6288_wire_96_31,
c6288_wire_96_32,
c6288_wire_96_33,
c6288_wire_96_34,
c6288_wire_96_35,
c6288_wire_96_36,
c6288_wire_96_37,
c6288_wire_96_38,
c6288_wire_96_39,
c6288_wire_96_40,
c6288_wire_96_41,
c6288_wire_96_42,
c6288_wire_96_43,
c6288_wire_96_44,
c6288_wire_96_45,
c6288_wire_96_46,
c6288_wire_99_0,
c6288_wire_99_1,
c6288_wire_99_2,
c6288_wire_99_3,
c6288_wire_99_4,
c6288_wire_99_5,
c6288_wire_99_6,
c6288_wire_99_7,
c6288_wire_99_8,
c6288_wire_99_9,
c6288_wire_99_10,
c6288_wire_99_11,
c6288_wire_99_12,
c6288_wire_99_13,
c6288_wire_99_14,
c6288_wire_99_15,
c6288_wire_99_16,
c6288_wire_99_17,
c6288_wire_99_18,
c6288_wire_99_19,
c6288_wire_99_20,
c6288_wire_99_21,
c6288_wire_99_22,
c6288_wire_99_23,
c6288_wire_99_24,
c6288_wire_99_25,
c6288_wire_99_26,
c6288_wire_99_27,
c6288_wire_99_28,
c6288_wire_99_29,
c6288_wire_99_30,
c6288_wire_99_31,
c6288_wire_99_32,
c6288_wire_99_33,
c6288_wire_99_34,
c6288_wire_99_35,
c6288_wire_99_36,
c6288_wire_99_37,
c6288_wire_99_38,
c6288_wire_99_39,
c6288_wire_99_40,
c6288_wire_99_41,
c6288_wire_99_42,
c6288_wire_99_43,
c6288_wire_99_44,
c6288_wire_99_45,
c6288_wire_99_46,
c6288_wire_102_0,
c6288_wire_102_1,
c6288_wire_102_2,
c6288_wire_102_3,
c6288_wire_102_4,
c6288_wire_102_5,
c6288_wire_102_6,
c6288_wire_102_7,
c6288_wire_102_8,
c6288_wire_102_9,
c6288_wire_102_10,
c6288_wire_102_11,
c6288_wire_102_12,
c6288_wire_102_13,
c6288_wire_102_14,
c6288_wire_102_15,
c6288_wire_102_16,
c6288_wire_102_17,
c6288_wire_102_18,
c6288_wire_102_19,
c6288_wire_102_20,
c6288_wire_102_21,
c6288_wire_102_22,
c6288_wire_102_23,
c6288_wire_102_24,
c6288_wire_102_25,
c6288_wire_102_26,
c6288_wire_102_27,
c6288_wire_102_28,
c6288_wire_102_29,
c6288_wire_102_30,
c6288_wire_102_31,
c6288_wire_102_32,
c6288_wire_102_33,
c6288_wire_102_34,
c6288_wire_102_35,
c6288_wire_102_36,
c6288_wire_102_37,
c6288_wire_102_38,
c6288_wire_102_39,
c6288_wire_102_40,
c6288_wire_102_41,
c6288_wire_102_42,
c6288_wire_102_43,
c6288_wire_102_44,
c6288_wire_102_45,
c6288_wire_102_46,
c6288_wire_105_0,
c6288_wire_105_1,
c6288_wire_105_2,
c6288_wire_105_3,
c6288_wire_105_4,
c6288_wire_105_5,
c6288_wire_105_6,
c6288_wire_105_7,
c6288_wire_105_8,
c6288_wire_105_9,
c6288_wire_105_10,
c6288_wire_105_11,
c6288_wire_105_12,
c6288_wire_105_13,
c6288_wire_105_14,
c6288_wire_105_15,
c6288_wire_105_16,
c6288_wire_105_17,
c6288_wire_105_18,
c6288_wire_105_19,
c6288_wire_105_20,
c6288_wire_105_21,
c6288_wire_105_22,
c6288_wire_105_23,
c6288_wire_105_24,
c6288_wire_105_25,
c6288_wire_105_26,
c6288_wire_105_27,
c6288_wire_105_28,
c6288_wire_105_29,
c6288_wire_105_30,
c6288_wire_105_31,
c6288_wire_105_32,
c6288_wire_105_33,
c6288_wire_105_34,
c6288_wire_105_35,
c6288_wire_105_36,
c6288_wire_105_37,
c6288_wire_105_38,
c6288_wire_105_39,
c6288_wire_105_40,
c6288_wire_105_41,
c6288_wire_105_42,
c6288_wire_105_43,
c6288_wire_105_44,
c6288_wire_105_45,
c6288_wire_105_46,
c6288_wire_108_0,
c6288_wire_108_1,
c6288_wire_108_2,
c6288_wire_108_3,
c6288_wire_108_4,
c6288_wire_108_5,
c6288_wire_108_6,
c6288_wire_108_7,
c6288_wire_108_8,
c6288_wire_108_9,
c6288_wire_108_10,
c6288_wire_108_11,
c6288_wire_108_12,
c6288_wire_108_13,
c6288_wire_108_14,
c6288_wire_108_15,
c6288_wire_108_16,
c6288_wire_108_17,
c6288_wire_108_18,
c6288_wire_108_19,
c6288_wire_108_20,
c6288_wire_108_21,
c6288_wire_108_22,
c6288_wire_108_23,
c6288_wire_108_24,
c6288_wire_108_25,
c6288_wire_108_26,
c6288_wire_108_27,
c6288_wire_108_28,
c6288_wire_108_29,
c6288_wire_108_30,
c6288_wire_108_31,
c6288_wire_108_32,
c6288_wire_108_33,
c6288_wire_108_34,
c6288_wire_108_35,
c6288_wire_108_36,
c6288_wire_108_37,
c6288_wire_108_38,
c6288_wire_108_39,
c6288_wire_108_40,
c6288_wire_108_41,
c6288_wire_108_42,
c6288_wire_108_43,
c6288_wire_108_44,
c6288_wire_108_45,
c6288_wire_108_46,
c6288_wire_111_0,
c6288_wire_111_1,
c6288_wire_111_2,
c6288_wire_111_3,
c6288_wire_111_4,
c6288_wire_111_5,
c6288_wire_111_6,
c6288_wire_111_7,
c6288_wire_111_8,
c6288_wire_111_9,
c6288_wire_111_10,
c6288_wire_111_11,
c6288_wire_111_12,
c6288_wire_111_13,
c6288_wire_111_14,
c6288_wire_111_15,
c6288_wire_111_16,
c6288_wire_111_17,
c6288_wire_111_18,
c6288_wire_111_19,
c6288_wire_111_20,
c6288_wire_111_21,
c6288_wire_111_22,
c6288_wire_111_23,
c6288_wire_111_24,
c6288_wire_111_25,
c6288_wire_111_26,
c6288_wire_111_27,
c6288_wire_111_28,
c6288_wire_111_29,
c6288_wire_111_30,
c6288_wire_111_31,
c6288_wire_111_32,
c6288_wire_111_33,
c6288_wire_111_34,
c6288_wire_111_35,
c6288_wire_111_36,
c6288_wire_111_37,
c6288_wire_111_38,
c6288_wire_111_39,
c6288_wire_111_40,
c6288_wire_111_41,
c6288_wire_111_42,
c6288_wire_111_43,
c6288_wire_111_44,
c6288_wire_111_45,
c6288_wire_111_46,
c6288_wire_114_0,
c6288_wire_114_1,
c6288_wire_114_2,
c6288_wire_114_3,
c6288_wire_114_4,
c6288_wire_114_5,
c6288_wire_114_6,
c6288_wire_114_7,
c6288_wire_114_8,
c6288_wire_114_9,
c6288_wire_114_10,
c6288_wire_114_11,
c6288_wire_114_12,
c6288_wire_114_13,
c6288_wire_114_14,
c6288_wire_114_15,
c6288_wire_114_16,
c6288_wire_114_17,
c6288_wire_114_18,
c6288_wire_114_19,
c6288_wire_114_20,
c6288_wire_114_21,
c6288_wire_114_22,
c6288_wire_114_23,
c6288_wire_114_24,
c6288_wire_114_25,
c6288_wire_114_26,
c6288_wire_114_27,
c6288_wire_114_28,
c6288_wire_114_29,
c6288_wire_114_30,
c6288_wire_114_31,
c6288_wire_114_32,
c6288_wire_114_33,
c6288_wire_114_34,
c6288_wire_114_35,
c6288_wire_114_36,
c6288_wire_114_37,
c6288_wire_114_38,
c6288_wire_114_39,
c6288_wire_114_40,
c6288_wire_114_41,
c6288_wire_114_42,
c6288_wire_114_43,
c6288_wire_114_44,
c6288_wire_114_45,
c6288_wire_114_46,
c6288_wire_42_0,
c6288_wire_42_1,
c6288_wire_42_2,
c6288_wire_42_3,
c6288_wire_42_4,
c6288_wire_42_5,
c6288_wire_42_6,
c6288_wire_42_7,
c6288_wire_42_8,
c6288_wire_42_9,
c6288_wire_42_10,
c6288_wire_42_11,
c6288_wire_42_12,
c6288_wire_42_13,
c6288_wire_42_14,
c6288_wire_42_15,
c6288_wire_42_16,
c6288_wire_42_17,
c6288_wire_42_18,
c6288_wire_42_19,
c6288_wire_42_20,
c6288_wire_42_21,
c6288_wire_42_22,
c6288_wire_42_23,
c6288_wire_42_24,
c6288_wire_42_25,
c6288_wire_42_26,
c6288_wire_42_27,
c6288_wire_42_28,
c6288_wire_42_29,
c6288_wire_42_30,
c6288_wire_42_31,
c6288_wire_42_32,
c6288_wire_42_33,
c6288_wire_42_34,
c6288_wire_42_35,
c6288_wire_42_36,
c6288_wire_42_37,
c6288_wire_42_38,
c6288_wire_42_39,
c6288_wire_42_40,
c6288_wire_42_41,
c6288_wire_42_42,
c6288_wire_42_43,
c6288_wire_42_44,
c6288_wire_42_45,
c6288_wire_117_0,
c6288_wire_117_1,
c6288_wire_117_2,
c6288_wire_117_3,
c6288_wire_117_4,
c6288_wire_117_5,
c6288_wire_117_6,
c6288_wire_117_7,
c6288_wire_117_8,
c6288_wire_117_9,
c6288_wire_117_10,
c6288_wire_117_11,
c6288_wire_117_12,
c6288_wire_117_13,
c6288_wire_117_14,
c6288_wire_117_15,
c6288_wire_117_16,
c6288_wire_117_17,
c6288_wire_117_18,
c6288_wire_117_19,
c6288_wire_117_20,
c6288_wire_117_21,
c6288_wire_117_22,
c6288_wire_117_23,
c6288_wire_117_24,
c6288_wire_117_25,
c6288_wire_117_26,
c6288_wire_117_27,
c6288_wire_117_28,
c6288_wire_117_29,
c6288_wire_117_30,
c6288_wire_117_31,
c6288_wire_117_32,
c6288_wire_117_33,
c6288_wire_117_34,
c6288_wire_117_35,
c6288_wire_117_36,
c6288_wire_117_37,
c6288_wire_117_38,
c6288_wire_117_39,
c6288_wire_117_40,
c6288_wire_117_41,
c6288_wire_117_42,
c6288_wire_117_43,
c6288_wire_117_44,
c6288_wire_117_45,
c6288_wire_117_46,
c6288_wire_47_0,
c6288_wire_47_1,
c6288_wire_47_2,
c6288_wire_47_3,
c6288_wire_47_4,
c6288_wire_47_5,
c6288_wire_47_6,
c6288_wire_47_7,
c6288_wire_47_8,
c6288_wire_47_9,
c6288_wire_47_10,
c6288_wire_47_11,
c6288_wire_47_12,
c6288_wire_47_13,
c6288_wire_47_14,
c6288_wire_47_15,
c6288_wire_47_16,
c6288_wire_47_17,
c6288_wire_47_18,
c6288_wire_47_19,
c6288_wire_47_20,
c6288_wire_47_21,
c6288_wire_47_22,
c6288_wire_47_23,
c6288_wire_47_24,
c6288_wire_47_25,
c6288_wire_47_26,
c6288_wire_47_27,
c6288_wire_47_28,
c6288_wire_47_29,
c6288_wire_47_30,
c6288_wire_47_31,
c6288_wire_47_32,
c6288_wire_47_33,
c6288_wire_47_34,
c6288_wire_47_35,
c6288_wire_47_36,
c6288_wire_47_37,
c6288_wire_47_38,
c6288_wire_47_39,
c6288_wire_47_40,
c6288_wire_47_41,
c6288_wire_47_42,
c6288_wire_47_43,
c6288_wire_47_44,
c6288_wire_47_45,
c6288_wire_52_0,
c6288_wire_52_1,
c6288_wire_52_2,
c6288_wire_52_3,
c6288_wire_52_4,
c6288_wire_52_5,
c6288_wire_52_6,
c6288_wire_52_7,
c6288_wire_52_8,
c6288_wire_52_9,
c6288_wire_52_10,
c6288_wire_52_11,
c6288_wire_52_12,
c6288_wire_52_13,
c6288_wire_52_14,
c6288_wire_52_15,
c6288_wire_52_16,
c6288_wire_52_17,
c6288_wire_52_18,
c6288_wire_52_19,
c6288_wire_52_20,
c6288_wire_52_21,
c6288_wire_52_22,
c6288_wire_52_23,
c6288_wire_52_24,
c6288_wire_52_25,
c6288_wire_52_26,
c6288_wire_52_27,
c6288_wire_52_28,
c6288_wire_52_29,
c6288_wire_52_30,
c6288_wire_52_31,
c6288_wire_52_32,
c6288_wire_52_33,
c6288_wire_52_34,
c6288_wire_52_35,
c6288_wire_52_36,
c6288_wire_52_37,
c6288_wire_52_38,
c6288_wire_52_39,
c6288_wire_52_40,
c6288_wire_52_41,
c6288_wire_52_42,
c6288_wire_52_43,
c6288_wire_52_44,
c6288_wire_52_45,
in256_net_0,
in239_net_0,
in222_net_0,
in205_net_0,
in188_net_0,
in171_net_0,
in154_net_0,
in137_net_0,
in120_net_0,
in103_net_0,
in86_net_0,
in69_net_0,
in52_net_0,
in35_net_0,
in18_net_0,
in1_net_0,
in528_net_0,
in511_net_0,
in494_net_0,
in477_net_0,
in460_net_0,
in443_net_0,
in426_net_0,
in409_net_0,
in392_net_0,
in375_net_0,
in358_net_0,
in341_net_0,
in324_net_0,
in307_net_0,
in290_net_0,
in273_net_0,
out6287_net_0,
out6288_net_0,
out6280_net_0,
out6270_net_0,
out6260_net_0,
out6250_net_0,
out6240_net_0,
out6230_net_0,
out6220_net_0,
out6210_net_0,
out6200_net_0,
out6190_net_0,
out6180_net_0,
out6170_net_0,
out6160_net_0,
out6150_net_0,
out6123_net_0,
out5971_net_0,
out5672_net_0,
out5308_net_0,
out4946_net_0,
out4591_net_0,
out4241_net_0,
out3895_net_0,
out3552_net_0,
out3211_net_0,
out2877_net_0,
out2548_net_0,
out2223_net_0,
out1901_net_0,
out1581_net_0,
out545_net_0;

pin #(32) pin_0 ({in256, in239, in222, in205, in188, in171, in154, in137, in120, in103, in86, in69, in52, in35, in18, in1, in528, in511, in494, in477, in460, in443, in426, in409, in392, in375, in358, in341, in324, in307, in290, in273}, {in256_net_0, in239_net_0, in222_net_0, in205_net_0, in188_net_0, in171_net_0, in154_net_0, in137_net_0, in120_net_0, in103_net_0, in86_net_0, in69_net_0, in52_net_0, in35_net_0, in18_net_0, in1_net_0, in528_net_0, in511_net_0, in494_net_0, in477_net_0, in460_net_0, in443_net_0, in426_net_0, in409_net_0, in392_net_0, in375_net_0, in358_net_0, in341_net_0, in324_net_0, in307_net_0, in290_net_0, in273_net_0});

pout #(32) pout_0 ({out6287_net_0, out6288_net_0, out6280_net_0, out6270_net_0, out6260_net_0, out6250_net_0, out6240_net_0, out6230_net_0, out6220_net_0, out6210_net_0, out6200_net_0, out6190_net_0, out6180_net_0, out6170_net_0, out6160_net_0, out6150_net_0, out6123_net_0, out5971_net_0, out5672_net_0, out5308_net_0, out4946_net_0, out4591_net_0, out4241_net_0, out3895_net_0, out3552_net_0, out3211_net_0, out2877_net_0, out2548_net_0, out2223_net_0, out1901_net_0, out1581_net_0, out545_net_0}, {out6287, out6288, out6280, out6270, out6260, out6250, out6240, out6230, out6220, out6210, out6200, out6190, out6180, out6170, out6160, out6150, out6123, out5971, out5672, out5308, out4946, out4591, out4241, out3895, out3552, out3211, out2877, out2548, out2223, out1901, out1581, out545});

fanout_n #(3, 0, 0) FANOUT_1 (c6288_wire_1, {c6288_wire_1_0, c6288_wire_1_1, c6288_wire_1_2});
fanout_n #(3, 0, 0) FANOUT_2 (c6288_wire_4, {c6288_wire_4_0, c6288_wire_4_1, c6288_wire_4_2});
fanout_n #(3, 0, 0) FANOUT_3 (c6288_wire_9, {c6288_wire_9_0, c6288_wire_9_1, c6288_wire_9_2});
fanout_n #(3, 0, 0) FANOUT_4 (c6288_wire_11, {c6288_wire_11_0, c6288_wire_11_1, c6288_wire_11_2});
fanout_n #(3, 0, 0) FANOUT_5 (c6288_wire_14, {c6288_wire_14_0, c6288_wire_14_1, c6288_wire_14_2});
fanout_n #(3, 0, 0) FANOUT_6 (c6288_wire_16, {c6288_wire_16_0, c6288_wire_16_1, c6288_wire_16_2});
fanout_n #(3, 0, 0) FANOUT_7 (c6288_wire_19, {c6288_wire_19_0, c6288_wire_19_1, c6288_wire_19_2});
fanout_n #(3, 0, 0) FANOUT_8 (c6288_wire_21, {c6288_wire_21_0, c6288_wire_21_1, c6288_wire_21_2});
fanout_n #(3, 0, 0) FANOUT_9 (c6288_wire_24, {c6288_wire_24_0, c6288_wire_24_1, c6288_wire_24_2});
fanout_n #(2, 0, 0) FANOUT_10 (c6288_wire_26, {c6288_wire_26_0, c6288_wire_26_1});
fanout_n #(3, 0, 0) FANOUT_11 (c6288_wire_29, {c6288_wire_29_0, c6288_wire_29_1, c6288_wire_29_2});
fanout_n #(3, 0, 0) FANOUT_12 (c6288_wire_31, {c6288_wire_31_0, c6288_wire_31_1, c6288_wire_31_2});
fanout_n #(3, 0, 0) FANOUT_13 (c6288_wire_36, {c6288_wire_36_0, c6288_wire_36_1, c6288_wire_36_2});
fanout_n #(3, 0, 0) FANOUT_14 (c6288_wire_38, {c6288_wire_38_0, c6288_wire_38_1, c6288_wire_38_2});
fanout_n #(3, 0, 0) FANOUT_15 (c6288_wire_41, {c6288_wire_41_0, c6288_wire_41_1, c6288_wire_41_2});
fanout_n #(3, 0, 0) FANOUT_16 (c6288_wire_43, {c6288_wire_43_0, c6288_wire_43_1, c6288_wire_43_2});
fanout_n #(3, 0, 0) FANOUT_17 (c6288_wire_46, {c6288_wire_46_0, c6288_wire_46_1, c6288_wire_46_2});
fanout_n #(3, 0, 0) FANOUT_18 (c6288_wire_48, {c6288_wire_48_0, c6288_wire_48_1, c6288_wire_48_2});
fanout_n #(3, 0, 0) FANOUT_19 (c6288_wire_51, {c6288_wire_51_0, c6288_wire_51_1, c6288_wire_51_2});
fanout_n #(3, 0, 0) FANOUT_20 (c6288_wire_53, {c6288_wire_53_0, c6288_wire_53_1, c6288_wire_53_2});
fanout_n #(3, 0, 0) FANOUT_21 (c6288_wire_56, {c6288_wire_56_0, c6288_wire_56_1, c6288_wire_56_2});
fanout_n #(3, 0, 0) FANOUT_22 (c6288_wire_58, {c6288_wire_58_0, c6288_wire_58_1, c6288_wire_58_2});
fanout_n #(3, 0, 0) FANOUT_23 (c6288_wire_61, {c6288_wire_61_0, c6288_wire_61_1, c6288_wire_61_2});
fanout_n #(3, 0, 0) FANOUT_24 (c6288_wire_63, {c6288_wire_63_0, c6288_wire_63_1, c6288_wire_63_2});
fanout_n #(3, 0, 0) FANOUT_25 (c6288_wire_66, {c6288_wire_66_0, c6288_wire_66_1, c6288_wire_66_2});
fanout_n #(3, 0, 0) FANOUT_26 (c6288_wire_68, {c6288_wire_68_0, c6288_wire_68_1, c6288_wire_68_2});
fanout_n #(3, 0, 0) FANOUT_27 (c6288_wire_71, {c6288_wire_71_0, c6288_wire_71_1, c6288_wire_71_2});
fanout_n #(3, 0, 0) FANOUT_28 (c6288_wire_72, {c6288_wire_72_0, c6288_wire_72_1, c6288_wire_72_2});
fanout_n #(3, 0, 0) FANOUT_29 (c6288_wire_327, {c6288_wire_327_0, c6288_wire_327_1, c6288_wire_327_2});
fanout_n #(3, 0, 0) FANOUT_30 (c6288_wire_748, {c6288_wire_748_0, c6288_wire_748_1, c6288_wire_748_2});
fanout_n #(2, 0, 0) FANOUT_31 (c6288_wire_749, {c6288_wire_749_0, c6288_wire_749_1});
fanout_n #(3, 0, 0) FANOUT_32 (c6288_wire_757, {c6288_wire_757_0, c6288_wire_757_1, c6288_wire_757_2});
fanout_n #(2, 0, 0) FANOUT_33 (c6288_wire_758, {c6288_wire_758_0, c6288_wire_758_1});
fanout_n #(3, 0, 0) FANOUT_34 (c6288_wire_763, {c6288_wire_763_0, c6288_wire_763_1, c6288_wire_763_2});
fanout_n #(2, 0, 0) FANOUT_35 (c6288_wire_764, {c6288_wire_764_0, c6288_wire_764_1});
fanout_n #(3, 0, 0) FANOUT_36 (c6288_wire_769, {c6288_wire_769_0, c6288_wire_769_1, c6288_wire_769_2});
fanout_n #(2, 0, 0) FANOUT_37 (c6288_wire_770, {c6288_wire_770_0, c6288_wire_770_1});
fanout_n #(2, 0, 0) FANOUT_38 (c6288_wire_776, {c6288_wire_776_0, c6288_wire_776_1});
fanout_n #(2, 0, 0) FANOUT_39 (c6288_wire_780, {c6288_wire_780_0, c6288_wire_780_1});
fanout_n #(3, 0, 0) FANOUT_40 (c6288_wire_784, {c6288_wire_784_0, c6288_wire_784_1, c6288_wire_784_2});
fanout_n #(2, 0, 0) FANOUT_41 (c6288_wire_785, {c6288_wire_785_0, c6288_wire_785_1});
fanout_n #(3, 0, 0) FANOUT_42 (c6288_wire_791, {c6288_wire_791_0, c6288_wire_791_1, c6288_wire_791_2});
fanout_n #(2, 0, 0) FANOUT_43 (c6288_wire_792, {c6288_wire_792_0, c6288_wire_792_1});
fanout_n #(3, 0, 0) FANOUT_44 (c6288_wire_797, {c6288_wire_797_0, c6288_wire_797_1, c6288_wire_797_2});
fanout_n #(2, 0, 0) FANOUT_45 (c6288_wire_798, {c6288_wire_798_0, c6288_wire_798_1});
fanout_n #(3, 0, 0) FANOUT_46 (c6288_wire_803, {c6288_wire_803_0, c6288_wire_803_1, c6288_wire_803_2});
fanout_n #(2, 0, 0) FANOUT_47 (c6288_wire_804, {c6288_wire_804_0, c6288_wire_804_1});
fanout_n #(3, 0, 0) FANOUT_48 (c6288_wire_809, {c6288_wire_809_0, c6288_wire_809_1, c6288_wire_809_2});
fanout_n #(2, 0, 0) FANOUT_49 (c6288_wire_810, {c6288_wire_810_0, c6288_wire_810_1});
fanout_n #(3, 0, 0) FANOUT_50 (c6288_wire_815, {c6288_wire_815_0, c6288_wire_815_1, c6288_wire_815_2});
fanout_n #(2, 0, 0) FANOUT_51 (c6288_wire_816, {c6288_wire_816_0, c6288_wire_816_1});
fanout_n #(3, 0, 0) FANOUT_52 (c6288_wire_821, {c6288_wire_821_0, c6288_wire_821_1, c6288_wire_821_2});
fanout_n #(2, 0, 0) FANOUT_53 (c6288_wire_822, {c6288_wire_822_0, c6288_wire_822_1});
fanout_n #(3, 0, 0) FANOUT_54 (c6288_wire_827, {c6288_wire_827_0, c6288_wire_827_1, c6288_wire_827_2});
fanout_n #(2, 0, 0) FANOUT_55 (c6288_wire_828, {c6288_wire_828_0, c6288_wire_828_1});
fanout_n #(3, 0, 0) FANOUT_56 (c6288_wire_833, {c6288_wire_833_0, c6288_wire_833_1, c6288_wire_833_2});
fanout_n #(2, 0, 0) FANOUT_57 (c6288_wire_754, {c6288_wire_754_0, c6288_wire_754_1});
fanout_n #(3, 0, 0) FANOUT_58 (c6288_wire_140, {c6288_wire_140_0, c6288_wire_140_1, c6288_wire_140_2});
fanout_n #(2, 0, 0) FANOUT_59 (c6288_wire_839, {c6288_wire_839_0, c6288_wire_839_1});
fanout_n #(3, 0, 0) FANOUT_60 (c6288_wire_138, {c6288_wire_138_0, c6288_wire_138_1, c6288_wire_138_2});
fanout_n #(2, 0, 0) FANOUT_61 (c6288_wire_847, {c6288_wire_847_0, c6288_wire_847_1});
fanout_n #(3, 0, 0) FANOUT_62 (c6288_wire_136, {c6288_wire_136_0, c6288_wire_136_1, c6288_wire_136_2});
fanout_n #(2, 0, 0) FANOUT_63 (c6288_wire_852, {c6288_wire_852_0, c6288_wire_852_1});
fanout_n #(3, 0, 0) FANOUT_64 (c6288_wire_134, {c6288_wire_134_0, c6288_wire_134_1, c6288_wire_134_2});
fanout_n #(2, 0, 0) FANOUT_65 (c6288_wire_857, {c6288_wire_857_0, c6288_wire_857_1});
fanout_n #(3, 0, 0) FANOUT_66 (c6288_wire_862, {c6288_wire_862_0, c6288_wire_862_1, c6288_wire_862_2});
fanout_n #(2, 0, 0) FANOUT_67 (c6288_wire_863, {c6288_wire_863_0, c6288_wire_863_1});
fanout_n #(3, 0, 0) FANOUT_68 (c6288_wire_869, {c6288_wire_869_0, c6288_wire_869_1, c6288_wire_869_2});
fanout_n #(3, 0, 0) FANOUT_69 (c6288_wire_158, {c6288_wire_158_0, c6288_wire_158_1, c6288_wire_158_2});
fanout_n #(2, 0, 0) FANOUT_70 (c6288_wire_874, {c6288_wire_874_0, c6288_wire_874_1});
fanout_n #(3, 0, 0) FANOUT_71 (c6288_wire_156, {c6288_wire_156_0, c6288_wire_156_1, c6288_wire_156_2});
fanout_n #(2, 0, 0) FANOUT_72 (c6288_wire_880, {c6288_wire_880_0, c6288_wire_880_1});
fanout_n #(3, 0, 0) FANOUT_73 (c6288_wire_154, {c6288_wire_154_0, c6288_wire_154_1, c6288_wire_154_2});
fanout_n #(2, 0, 0) FANOUT_74 (c6288_wire_885, {c6288_wire_885_0, c6288_wire_885_1});
fanout_n #(3, 0, 0) FANOUT_75 (c6288_wire_152, {c6288_wire_152_0, c6288_wire_152_1, c6288_wire_152_2});
fanout_n #(2, 0, 0) FANOUT_76 (c6288_wire_890, {c6288_wire_890_0, c6288_wire_890_1});
fanout_n #(3, 0, 0) FANOUT_77 (c6288_wire_150, {c6288_wire_150_0, c6288_wire_150_1, c6288_wire_150_2});
fanout_n #(2, 0, 0) FANOUT_78 (c6288_wire_895, {c6288_wire_895_0, c6288_wire_895_1});
fanout_n #(3, 0, 0) FANOUT_79 (c6288_wire_148, {c6288_wire_148_0, c6288_wire_148_1, c6288_wire_148_2});
fanout_n #(2, 0, 0) FANOUT_80 (c6288_wire_900, {c6288_wire_900_0, c6288_wire_900_1});
fanout_n #(3, 0, 0) FANOUT_81 (c6288_wire_146, {c6288_wire_146_0, c6288_wire_146_1, c6288_wire_146_2});
fanout_n #(2, 0, 0) FANOUT_82 (c6288_wire_905, {c6288_wire_905_0, c6288_wire_905_1});
fanout_n #(3, 0, 0) FANOUT_83 (c6288_wire_144, {c6288_wire_144_0, c6288_wire_144_1, c6288_wire_144_2});
fanout_n #(2, 0, 0) FANOUT_84 (c6288_wire_910, {c6288_wire_910_0, c6288_wire_910_1});
fanout_n #(3, 0, 0) FANOUT_85 (c6288_wire_142, {c6288_wire_142_0, c6288_wire_142_1, c6288_wire_142_2});
fanout_n #(2, 0, 0) FANOUT_86 (c6288_wire_844, {c6288_wire_844_0, c6288_wire_844_1});
fanout_n #(3, 0, 0) FANOUT_87 (c6288_wire_182, {c6288_wire_182_0, c6288_wire_182_1, c6288_wire_182_2});
fanout_n #(2, 0, 0) FANOUT_88 (c6288_wire_920, {c6288_wire_920_0, c6288_wire_920_1});
fanout_n #(3, 0, 0) FANOUT_89 (c6288_wire_180, {c6288_wire_180_0, c6288_wire_180_1, c6288_wire_180_2});
fanout_n #(2, 0, 0) FANOUT_90 (c6288_wire_928, {c6288_wire_928_0, c6288_wire_928_1});
fanout_n #(3, 0, 0) FANOUT_91 (c6288_wire_178, {c6288_wire_178_0, c6288_wire_178_1, c6288_wire_178_2});
fanout_n #(2, 0, 0) FANOUT_92 (c6288_wire_933, {c6288_wire_933_0, c6288_wire_933_1});
fanout_n #(3, 0, 0) FANOUT_93 (c6288_wire_176, {c6288_wire_176_0, c6288_wire_176_1, c6288_wire_176_2});
fanout_n #(2, 0, 0) FANOUT_94 (c6288_wire_938, {c6288_wire_938_0, c6288_wire_938_1});
fanout_n #(3, 0, 0) FANOUT_95 (c6288_wire_870, {c6288_wire_870_0, c6288_wire_870_1, c6288_wire_870_2});
fanout_n #(2, 0, 0) FANOUT_96 (c6288_wire_943, {c6288_wire_943_0, c6288_wire_943_1});
fanout_n #(3, 0, 0) FANOUT_97 (c6288_wire_949, {c6288_wire_949_0, c6288_wire_949_1, c6288_wire_949_2});
fanout_n #(3, 0, 0) FANOUT_98 (c6288_wire_200, {c6288_wire_200_0, c6288_wire_200_1, c6288_wire_200_2});
fanout_n #(2, 0, 0) FANOUT_99 (c6288_wire_952, {c6288_wire_952_0, c6288_wire_952_1});
fanout_n #(3, 0, 0) FANOUT_100 (c6288_wire_198, {c6288_wire_198_0, c6288_wire_198_1, c6288_wire_198_2});
fanout_n #(2, 0, 0) FANOUT_101 (c6288_wire_958, {c6288_wire_958_0, c6288_wire_958_1});
fanout_n #(3, 0, 0) FANOUT_102 (c6288_wire_196, {c6288_wire_196_0, c6288_wire_196_1, c6288_wire_196_2});
fanout_n #(2, 0, 0) FANOUT_103 (c6288_wire_963, {c6288_wire_963_0, c6288_wire_963_1});
fanout_n #(3, 0, 0) FANOUT_104 (c6288_wire_194, {c6288_wire_194_0, c6288_wire_194_1, c6288_wire_194_2});
fanout_n #(2, 0, 0) FANOUT_105 (c6288_wire_968, {c6288_wire_968_0, c6288_wire_968_1});
fanout_n #(3, 0, 0) FANOUT_106 (c6288_wire_192, {c6288_wire_192_0, c6288_wire_192_1, c6288_wire_192_2});
fanout_n #(2, 0, 0) FANOUT_107 (c6288_wire_973, {c6288_wire_973_0, c6288_wire_973_1});
fanout_n #(3, 0, 0) FANOUT_108 (c6288_wire_190, {c6288_wire_190_0, c6288_wire_190_1, c6288_wire_190_2});
fanout_n #(2, 0, 0) FANOUT_109 (c6288_wire_978, {c6288_wire_978_0, c6288_wire_978_1});
fanout_n #(3, 0, 0) FANOUT_110 (c6288_wire_188, {c6288_wire_188_0, c6288_wire_188_1, c6288_wire_188_2});
fanout_n #(2, 0, 0) FANOUT_111 (c6288_wire_983, {c6288_wire_983_0, c6288_wire_983_1});
fanout_n #(3, 0, 0) FANOUT_112 (c6288_wire_186, {c6288_wire_186_0, c6288_wire_186_1, c6288_wire_186_2});
fanout_n #(2, 0, 0) FANOUT_113 (c6288_wire_988, {c6288_wire_988_0, c6288_wire_988_1});
fanout_n #(3, 0, 0) FANOUT_114 (c6288_wire_184, {c6288_wire_184_0, c6288_wire_184_1, c6288_wire_184_2});
fanout_n #(2, 0, 0) FANOUT_115 (c6288_wire_925, {c6288_wire_925_0, c6288_wire_925_1});
fanout_n #(3, 0, 0) FANOUT_116 (c6288_wire_224, {c6288_wire_224_0, c6288_wire_224_1, c6288_wire_224_2});
fanout_n #(2, 0, 0) FANOUT_117 (c6288_wire_998, {c6288_wire_998_0, c6288_wire_998_1});
fanout_n #(3, 0, 0) FANOUT_118 (c6288_wire_222, {c6288_wire_222_0, c6288_wire_222_1, c6288_wire_222_2});
fanout_n #(2, 0, 0) FANOUT_119 (c6288_wire_1006, {c6288_wire_1006_0, c6288_wire_1006_1});
fanout_n #(3, 0, 0) FANOUT_120 (c6288_wire_220, {c6288_wire_220_0, c6288_wire_220_1, c6288_wire_220_2});
fanout_n #(2, 0, 0) FANOUT_121 (c6288_wire_1011, {c6288_wire_1011_0, c6288_wire_1011_1});
fanout_n #(3, 0, 0) FANOUT_122 (c6288_wire_218, {c6288_wire_218_0, c6288_wire_218_1, c6288_wire_218_2});
fanout_n #(2, 0, 0) FANOUT_123 (c6288_wire_1016, {c6288_wire_1016_0, c6288_wire_1016_1});
fanout_n #(3, 0, 0) FANOUT_124 (c6288_wire_950, {c6288_wire_950_0, c6288_wire_950_1, c6288_wire_950_2});
fanout_n #(2, 0, 0) FANOUT_125 (c6288_wire_1021, {c6288_wire_1021_0, c6288_wire_1021_1});
fanout_n #(3, 0, 0) FANOUT_126 (c6288_wire_1027, {c6288_wire_1027_0, c6288_wire_1027_1, c6288_wire_1027_2});
fanout_n #(3, 0, 0) FANOUT_127 (c6288_wire_242, {c6288_wire_242_0, c6288_wire_242_1, c6288_wire_242_2});
fanout_n #(2, 0, 0) FANOUT_128 (c6288_wire_1030, {c6288_wire_1030_0, c6288_wire_1030_1});
fanout_n #(3, 0, 0) FANOUT_129 (c6288_wire_240, {c6288_wire_240_0, c6288_wire_240_1, c6288_wire_240_2});
fanout_n #(2, 0, 0) FANOUT_130 (c6288_wire_1036, {c6288_wire_1036_0, c6288_wire_1036_1});
fanout_n #(3, 0, 0) FANOUT_131 (c6288_wire_238, {c6288_wire_238_0, c6288_wire_238_1, c6288_wire_238_2});
fanout_n #(2, 0, 0) FANOUT_132 (c6288_wire_1041, {c6288_wire_1041_0, c6288_wire_1041_1});
fanout_n #(3, 0, 0) FANOUT_133 (c6288_wire_236, {c6288_wire_236_0, c6288_wire_236_1, c6288_wire_236_2});
fanout_n #(2, 0, 0) FANOUT_134 (c6288_wire_1046, {c6288_wire_1046_0, c6288_wire_1046_1});
fanout_n #(3, 0, 0) FANOUT_135 (c6288_wire_234, {c6288_wire_234_0, c6288_wire_234_1, c6288_wire_234_2});
fanout_n #(2, 0, 0) FANOUT_136 (c6288_wire_1051, {c6288_wire_1051_0, c6288_wire_1051_1});
fanout_n #(3, 0, 0) FANOUT_137 (c6288_wire_232, {c6288_wire_232_0, c6288_wire_232_1, c6288_wire_232_2});
fanout_n #(2, 0, 0) FANOUT_138 (c6288_wire_1056, {c6288_wire_1056_0, c6288_wire_1056_1});
fanout_n #(3, 0, 0) FANOUT_139 (c6288_wire_230, {c6288_wire_230_0, c6288_wire_230_1, c6288_wire_230_2});
fanout_n #(2, 0, 0) FANOUT_140 (c6288_wire_1061, {c6288_wire_1061_0, c6288_wire_1061_1});
fanout_n #(3, 0, 0) FANOUT_141 (c6288_wire_228, {c6288_wire_228_0, c6288_wire_228_1, c6288_wire_228_2});
fanout_n #(2, 0, 0) FANOUT_142 (c6288_wire_1066, {c6288_wire_1066_0, c6288_wire_1066_1});
fanout_n #(3, 0, 0) FANOUT_143 (c6288_wire_226, {c6288_wire_226_0, c6288_wire_226_1, c6288_wire_226_2});
fanout_n #(2, 0, 0) FANOUT_144 (c6288_wire_1003, {c6288_wire_1003_0, c6288_wire_1003_1});
fanout_n #(3, 0, 0) FANOUT_145 (c6288_wire_286, {c6288_wire_286_0, c6288_wire_286_1, c6288_wire_286_2});
fanout_n #(3, 0, 0) FANOUT_146 (c6288_wire_266, {c6288_wire_266_0, c6288_wire_266_1, c6288_wire_266_2});
fanout_n #(2, 0, 0) FANOUT_147 (c6288_wire_1074, {c6288_wire_1074_0, c6288_wire_1074_1});
fanout_n #(3, 0, 0) FANOUT_148 (c6288_wire_264, {c6288_wire_264_0, c6288_wire_264_1, c6288_wire_264_2});
fanout_n #(2, 0, 0) FANOUT_149 (c6288_wire_1082, {c6288_wire_1082_0, c6288_wire_1082_1});
fanout_n #(3, 0, 0) FANOUT_150 (c6288_wire_262, {c6288_wire_262_0, c6288_wire_262_1, c6288_wire_262_2});
fanout_n #(2, 0, 0) FANOUT_151 (c6288_wire_1087, {c6288_wire_1087_0, c6288_wire_1087_1});
fanout_n #(3, 0, 0) FANOUT_152 (c6288_wire_260, {c6288_wire_260_0, c6288_wire_260_1, c6288_wire_260_2});
fanout_n #(2, 0, 0) FANOUT_153 (c6288_wire_1092, {c6288_wire_1092_0, c6288_wire_1092_1});
fanout_n #(3, 0, 0) FANOUT_154 (c6288_wire_1028, {c6288_wire_1028_0, c6288_wire_1028_1, c6288_wire_1028_2});
fanout_n #(2, 0, 0) FANOUT_155 (c6288_wire_1097, {c6288_wire_1097_0, c6288_wire_1097_1});
fanout_n #(4, 0, 0) FANOUT_156 (c6288_wire_1103, {c6288_wire_1103_0, c6288_wire_1103_1, c6288_wire_1103_2, c6288_wire_1103_3});
fanout_n #(3, 0, 0) FANOUT_157 (c6288_wire_1108, {c6288_wire_1108_0, c6288_wire_1108_1, c6288_wire_1108_2});
fanout_n #(3, 0, 0) FANOUT_158 (c6288_wire_282, {c6288_wire_282_0, c6288_wire_282_1, c6288_wire_282_2});
fanout_n #(2, 0, 0) FANOUT_159 (c6288_wire_1115, {c6288_wire_1115_0, c6288_wire_1115_1});
fanout_n #(3, 0, 0) FANOUT_160 (c6288_wire_280, {c6288_wire_280_0, c6288_wire_280_1, c6288_wire_280_2});
fanout_n #(2, 0, 0) FANOUT_161 (c6288_wire_1120, {c6288_wire_1120_0, c6288_wire_1120_1});
fanout_n #(3, 0, 0) FANOUT_162 (c6288_wire_278, {c6288_wire_278_0, c6288_wire_278_1, c6288_wire_278_2});
fanout_n #(2, 0, 0) FANOUT_163 (c6288_wire_1125, {c6288_wire_1125_0, c6288_wire_1125_1});
fanout_n #(3, 0, 0) FANOUT_164 (c6288_wire_276, {c6288_wire_276_0, c6288_wire_276_1, c6288_wire_276_2});
fanout_n #(2, 0, 0) FANOUT_165 (c6288_wire_1130, {c6288_wire_1130_0, c6288_wire_1130_1});
fanout_n #(3, 0, 0) FANOUT_166 (c6288_wire_274, {c6288_wire_274_0, c6288_wire_274_1, c6288_wire_274_2});
fanout_n #(2, 0, 0) FANOUT_167 (c6288_wire_1135, {c6288_wire_1135_0, c6288_wire_1135_1});
fanout_n #(3, 0, 0) FANOUT_168 (c6288_wire_272, {c6288_wire_272_0, c6288_wire_272_1, c6288_wire_272_2});
fanout_n #(2, 0, 0) FANOUT_169 (c6288_wire_1140, {c6288_wire_1140_0, c6288_wire_1140_1});
fanout_n #(3, 0, 0) FANOUT_170 (c6288_wire_270, {c6288_wire_270_0, c6288_wire_270_1, c6288_wire_270_2});
fanout_n #(2, 0, 0) FANOUT_171 (c6288_wire_1145, {c6288_wire_1145_0, c6288_wire_1145_1});
fanout_n #(3, 0, 0) FANOUT_172 (c6288_wire_268, {c6288_wire_268_0, c6288_wire_268_1, c6288_wire_268_2});
fanout_n #(2, 0, 0) FANOUT_173 (c6288_wire_1079, {c6288_wire_1079_0, c6288_wire_1079_1});
fanout_n #(3, 0, 0) FANOUT_174 (c6288_wire_1152, {c6288_wire_1152_0, c6288_wire_1152_1, c6288_wire_1152_2});
fanout_n #(3, 0, 0) FANOUT_175 (c6288_wire_1159, {c6288_wire_1159_0, c6288_wire_1159_1, c6288_wire_1159_2});
fanout_n #(3, 0, 0) FANOUT_176 (c6288_wire_1165, {c6288_wire_1165_0, c6288_wire_1165_1, c6288_wire_1165_2});
fanout_n #(3, 0, 0) FANOUT_177 (c6288_wire_1171, {c6288_wire_1171_0, c6288_wire_1171_1, c6288_wire_1171_2});
fanout_n #(4, 0, 0) FANOUT_178 (c6288_wire_1177, {c6288_wire_1177_0, c6288_wire_1177_1, c6288_wire_1177_2, c6288_wire_1177_3});
fanout_n #(3, 0, 0) FANOUT_179 (c6288_wire_1186, {c6288_wire_1186_0, c6288_wire_1186_1, c6288_wire_1186_2});
fanout_n #(3, 0, 0) FANOUT_180 (c6288_wire_1192, {c6288_wire_1192_0, c6288_wire_1192_1, c6288_wire_1192_2});
fanout_n #(3, 0, 0) FANOUT_181 (c6288_wire_1198, {c6288_wire_1198_0, c6288_wire_1198_1, c6288_wire_1198_2});
fanout_n #(3, 0, 0) FANOUT_182 (c6288_wire_1204, {c6288_wire_1204_0, c6288_wire_1204_1, c6288_wire_1204_2});
fanout_n #(3, 0, 0) FANOUT_183 (c6288_wire_1210, {c6288_wire_1210_0, c6288_wire_1210_1, c6288_wire_1210_2});
fanout_n #(3, 0, 0) FANOUT_184 (c6288_wire_1216, {c6288_wire_1216_0, c6288_wire_1216_1, c6288_wire_1216_2});
fanout_n #(3, 0, 0) FANOUT_185 (c6288_wire_1222, {c6288_wire_1222_0, c6288_wire_1222_1, c6288_wire_1222_2});
fanout_n #(3, 0, 0) FANOUT_186 (c6288_wire_1228, {c6288_wire_1228_0, c6288_wire_1228_1, c6288_wire_1228_2});
fanout_n #(3, 0, 0) FANOUT_187 (c6288_wire_382, {c6288_wire_382_0, c6288_wire_382_1, c6288_wire_382_2});
fanout_n #(2, 0, 0) FANOUT_188 (c6288_wire_1236, {c6288_wire_1236_0, c6288_wire_1236_1});
fanout_n #(3, 0, 0) FANOUT_189 (c6288_wire_380, {c6288_wire_380_0, c6288_wire_380_1, c6288_wire_380_2});
fanout_n #(2, 0, 0) FANOUT_190 (c6288_wire_1244, {c6288_wire_1244_0, c6288_wire_1244_1});
fanout_n #(3, 0, 0) FANOUT_191 (c6288_wire_378, {c6288_wire_378_0, c6288_wire_378_1, c6288_wire_378_2});
fanout_n #(2, 0, 0) FANOUT_192 (c6288_wire_1249, {c6288_wire_1249_0, c6288_wire_1249_1});
fanout_n #(3, 0, 0) FANOUT_193 (c6288_wire_376, {c6288_wire_376_0, c6288_wire_376_1, c6288_wire_376_2});
fanout_n #(2, 0, 0) FANOUT_194 (c6288_wire_1254, {c6288_wire_1254_0, c6288_wire_1254_1});
fanout_n #(2, 0, 0) FANOUT_195 (c6288_wire_782, {c6288_wire_782_0, c6288_wire_782_1});
fanout_n #(2, 0, 0) FANOUT_196 (c6288_wire_1259, {c6288_wire_1259_0, c6288_wire_1259_1});
fanout_n #(3, 0, 0) FANOUT_197 (c6288_wire_1265, {c6288_wire_1265_0, c6288_wire_1265_1, c6288_wire_1265_2});
fanout_n #(3, 0, 0) FANOUT_198 (c6288_wire_400, {c6288_wire_400_0, c6288_wire_400_1, c6288_wire_400_2});
fanout_n #(2, 0, 0) FANOUT_199 (c6288_wire_1269, {c6288_wire_1269_0, c6288_wire_1269_1});
fanout_n #(3, 0, 0) FANOUT_200 (c6288_wire_398, {c6288_wire_398_0, c6288_wire_398_1, c6288_wire_398_2});
fanout_n #(2, 0, 0) FANOUT_201 (c6288_wire_1275, {c6288_wire_1275_0, c6288_wire_1275_1});
fanout_n #(3, 0, 0) FANOUT_202 (c6288_wire_396, {c6288_wire_396_0, c6288_wire_396_1, c6288_wire_396_2});
fanout_n #(2, 0, 0) FANOUT_203 (c6288_wire_1280, {c6288_wire_1280_0, c6288_wire_1280_1});
fanout_n #(3, 0, 0) FANOUT_204 (c6288_wire_394, {c6288_wire_394_0, c6288_wire_394_1, c6288_wire_394_2});
fanout_n #(2, 0, 0) FANOUT_205 (c6288_wire_1285, {c6288_wire_1285_0, c6288_wire_1285_1});
fanout_n #(3, 0, 0) FANOUT_206 (c6288_wire_392, {c6288_wire_392_0, c6288_wire_392_1, c6288_wire_392_2});
fanout_n #(2, 0, 0) FANOUT_207 (c6288_wire_1290, {c6288_wire_1290_0, c6288_wire_1290_1});
fanout_n #(3, 0, 0) FANOUT_208 (c6288_wire_390, {c6288_wire_390_0, c6288_wire_390_1, c6288_wire_390_2});
fanout_n #(2, 0, 0) FANOUT_209 (c6288_wire_1295, {c6288_wire_1295_0, c6288_wire_1295_1});
fanout_n #(3, 0, 0) FANOUT_210 (c6288_wire_388, {c6288_wire_388_0, c6288_wire_388_1, c6288_wire_388_2});
fanout_n #(2, 0, 0) FANOUT_211 (c6288_wire_1300, {c6288_wire_1300_0, c6288_wire_1300_1});
fanout_n #(3, 0, 0) FANOUT_212 (c6288_wire_386, {c6288_wire_386_0, c6288_wire_386_1, c6288_wire_386_2});
fanout_n #(2, 0, 0) FANOUT_213 (c6288_wire_1305, {c6288_wire_1305_0, c6288_wire_1305_1});
fanout_n #(3, 0, 0) FANOUT_214 (c6288_wire_384, {c6288_wire_384_0, c6288_wire_384_1, c6288_wire_384_2});
fanout_n #(2, 0, 0) FANOUT_215 (c6288_wire_1241, {c6288_wire_1241_0, c6288_wire_1241_1});
fanout_n #(3, 0, 0) FANOUT_216 (c6288_wire_424, {c6288_wire_424_0, c6288_wire_424_1, c6288_wire_424_2});
fanout_n #(2, 0, 0) FANOUT_217 (c6288_wire_1315, {c6288_wire_1315_0, c6288_wire_1315_1});
fanout_n #(3, 0, 0) FANOUT_218 (c6288_wire_422, {c6288_wire_422_0, c6288_wire_422_1, c6288_wire_422_2});
fanout_n #(2, 0, 0) FANOUT_219 (c6288_wire_1323, {c6288_wire_1323_0, c6288_wire_1323_1});
fanout_n #(3, 0, 0) FANOUT_220 (c6288_wire_420, {c6288_wire_420_0, c6288_wire_420_1, c6288_wire_420_2});
fanout_n #(2, 0, 0) FANOUT_221 (c6288_wire_1328, {c6288_wire_1328_0, c6288_wire_1328_1});
fanout_n #(3, 0, 0) FANOUT_222 (c6288_wire_418, {c6288_wire_418_0, c6288_wire_418_1, c6288_wire_418_2});
fanout_n #(2, 0, 0) FANOUT_223 (c6288_wire_1333, {c6288_wire_1333_0, c6288_wire_1333_1});
fanout_n #(3, 0, 0) FANOUT_224 (c6288_wire_1266, {c6288_wire_1266_0, c6288_wire_1266_1, c6288_wire_1266_2});
fanout_n #(2, 0, 0) FANOUT_225 (c6288_wire_1338, {c6288_wire_1338_0, c6288_wire_1338_1});
fanout_n #(3, 0, 0) FANOUT_226 (c6288_wire_1344, {c6288_wire_1344_0, c6288_wire_1344_1, c6288_wire_1344_2});
fanout_n #(3, 0, 0) FANOUT_227 (c6288_wire_442, {c6288_wire_442_0, c6288_wire_442_1, c6288_wire_442_2});
fanout_n #(2, 0, 0) FANOUT_228 (c6288_wire_1347, {c6288_wire_1347_0, c6288_wire_1347_1});
fanout_n #(3, 0, 0) FANOUT_229 (c6288_wire_440, {c6288_wire_440_0, c6288_wire_440_1, c6288_wire_440_2});
fanout_n #(2, 0, 0) FANOUT_230 (c6288_wire_1353, {c6288_wire_1353_0, c6288_wire_1353_1});
fanout_n #(3, 0, 0) FANOUT_231 (c6288_wire_438, {c6288_wire_438_0, c6288_wire_438_1, c6288_wire_438_2});
fanout_n #(2, 0, 0) FANOUT_232 (c6288_wire_1358, {c6288_wire_1358_0, c6288_wire_1358_1});
fanout_n #(3, 0, 0) FANOUT_233 (c6288_wire_436, {c6288_wire_436_0, c6288_wire_436_1, c6288_wire_436_2});
fanout_n #(2, 0, 0) FANOUT_234 (c6288_wire_1363, {c6288_wire_1363_0, c6288_wire_1363_1});
fanout_n #(3, 0, 0) FANOUT_235 (c6288_wire_434, {c6288_wire_434_0, c6288_wire_434_1, c6288_wire_434_2});
fanout_n #(2, 0, 0) FANOUT_236 (c6288_wire_1368, {c6288_wire_1368_0, c6288_wire_1368_1});
fanout_n #(3, 0, 0) FANOUT_237 (c6288_wire_432, {c6288_wire_432_0, c6288_wire_432_1, c6288_wire_432_2});
fanout_n #(2, 0, 0) FANOUT_238 (c6288_wire_1373, {c6288_wire_1373_0, c6288_wire_1373_1});
fanout_n #(3, 0, 0) FANOUT_239 (c6288_wire_430, {c6288_wire_430_0, c6288_wire_430_1, c6288_wire_430_2});
fanout_n #(2, 0, 0) FANOUT_240 (c6288_wire_1378, {c6288_wire_1378_0, c6288_wire_1378_1});
fanout_n #(3, 0, 0) FANOUT_241 (c6288_wire_428, {c6288_wire_428_0, c6288_wire_428_1, c6288_wire_428_2});
fanout_n #(2, 0, 0) FANOUT_242 (c6288_wire_1383, {c6288_wire_1383_0, c6288_wire_1383_1});
fanout_n #(3, 0, 0) FANOUT_243 (c6288_wire_426, {c6288_wire_426_0, c6288_wire_426_1, c6288_wire_426_2});
fanout_n #(2, 0, 0) FANOUT_244 (c6288_wire_1320, {c6288_wire_1320_0, c6288_wire_1320_1});
fanout_n #(3, 0, 0) FANOUT_245 (c6288_wire_466, {c6288_wire_466_0, c6288_wire_466_1, c6288_wire_466_2});
fanout_n #(2, 0, 0) FANOUT_246 (c6288_wire_1393, {c6288_wire_1393_0, c6288_wire_1393_1});
fanout_n #(3, 0, 0) FANOUT_247 (c6288_wire_464, {c6288_wire_464_0, c6288_wire_464_1, c6288_wire_464_2});
fanout_n #(2, 0, 0) FANOUT_248 (c6288_wire_1401, {c6288_wire_1401_0, c6288_wire_1401_1});
fanout_n #(3, 0, 0) FANOUT_249 (c6288_wire_462, {c6288_wire_462_0, c6288_wire_462_1, c6288_wire_462_2});
fanout_n #(2, 0, 0) FANOUT_250 (c6288_wire_1406, {c6288_wire_1406_0, c6288_wire_1406_1});
fanout_n #(3, 0, 0) FANOUT_251 (c6288_wire_460, {c6288_wire_460_0, c6288_wire_460_1, c6288_wire_460_2});
fanout_n #(2, 0, 0) FANOUT_252 (c6288_wire_1411, {c6288_wire_1411_0, c6288_wire_1411_1});
fanout_n #(3, 0, 0) FANOUT_253 (c6288_wire_1345, {c6288_wire_1345_0, c6288_wire_1345_1, c6288_wire_1345_2});
fanout_n #(2, 0, 0) FANOUT_254 (c6288_wire_1416, {c6288_wire_1416_0, c6288_wire_1416_1});
fanout_n #(3, 0, 0) FANOUT_255 (c6288_wire_1422, {c6288_wire_1422_0, c6288_wire_1422_1, c6288_wire_1422_2});
fanout_n #(3, 0, 0) FANOUT_256 (c6288_wire_484, {c6288_wire_484_0, c6288_wire_484_1, c6288_wire_484_2});
fanout_n #(2, 0, 0) FANOUT_257 (c6288_wire_1425, {c6288_wire_1425_0, c6288_wire_1425_1});
fanout_n #(3, 0, 0) FANOUT_258 (c6288_wire_482, {c6288_wire_482_0, c6288_wire_482_1, c6288_wire_482_2});
fanout_n #(2, 0, 0) FANOUT_259 (c6288_wire_1431, {c6288_wire_1431_0, c6288_wire_1431_1});
fanout_n #(3, 0, 0) FANOUT_260 (c6288_wire_480, {c6288_wire_480_0, c6288_wire_480_1, c6288_wire_480_2});
fanout_n #(2, 0, 0) FANOUT_261 (c6288_wire_1436, {c6288_wire_1436_0, c6288_wire_1436_1});
fanout_n #(3, 0, 0) FANOUT_262 (c6288_wire_478, {c6288_wire_478_0, c6288_wire_478_1, c6288_wire_478_2});
fanout_n #(2, 0, 0) FANOUT_263 (c6288_wire_1441, {c6288_wire_1441_0, c6288_wire_1441_1});
fanout_n #(3, 0, 0) FANOUT_264 (c6288_wire_476, {c6288_wire_476_0, c6288_wire_476_1, c6288_wire_476_2});
fanout_n #(2, 0, 0) FANOUT_265 (c6288_wire_1446, {c6288_wire_1446_0, c6288_wire_1446_1});
fanout_n #(3, 0, 0) FANOUT_266 (c6288_wire_474, {c6288_wire_474_0, c6288_wire_474_1, c6288_wire_474_2});
fanout_n #(2, 0, 0) FANOUT_267 (c6288_wire_1451, {c6288_wire_1451_0, c6288_wire_1451_1});
fanout_n #(3, 0, 0) FANOUT_268 (c6288_wire_472, {c6288_wire_472_0, c6288_wire_472_1, c6288_wire_472_2});
fanout_n #(2, 0, 0) FANOUT_269 (c6288_wire_1456, {c6288_wire_1456_0, c6288_wire_1456_1});
fanout_n #(3, 0, 0) FANOUT_270 (c6288_wire_470, {c6288_wire_470_0, c6288_wire_470_1, c6288_wire_470_2});
fanout_n #(2, 0, 0) FANOUT_271 (c6288_wire_1461, {c6288_wire_1461_0, c6288_wire_1461_1});
fanout_n #(3, 0, 0) FANOUT_272 (c6288_wire_468, {c6288_wire_468_0, c6288_wire_468_1, c6288_wire_468_2});
fanout_n #(2, 0, 0) FANOUT_273 (c6288_wire_1398, {c6288_wire_1398_0, c6288_wire_1398_1});
fanout_n #(3, 0, 0) FANOUT_274 (c6288_wire_508, {c6288_wire_508_0, c6288_wire_508_1, c6288_wire_508_2});
fanout_n #(2, 0, 0) FANOUT_275 (c6288_wire_1471, {c6288_wire_1471_0, c6288_wire_1471_1});
fanout_n #(3, 0, 0) FANOUT_276 (c6288_wire_506, {c6288_wire_506_0, c6288_wire_506_1, c6288_wire_506_2});
fanout_n #(2, 0, 0) FANOUT_277 (c6288_wire_1479, {c6288_wire_1479_0, c6288_wire_1479_1});
fanout_n #(3, 0, 0) FANOUT_278 (c6288_wire_504, {c6288_wire_504_0, c6288_wire_504_1, c6288_wire_504_2});
fanout_n #(2, 0, 0) FANOUT_279 (c6288_wire_1484, {c6288_wire_1484_0, c6288_wire_1484_1});
fanout_n #(3, 0, 0) FANOUT_280 (c6288_wire_502, {c6288_wire_502_0, c6288_wire_502_1, c6288_wire_502_2});
fanout_n #(2, 0, 0) FANOUT_281 (c6288_wire_1489, {c6288_wire_1489_0, c6288_wire_1489_1});
fanout_n #(3, 0, 0) FANOUT_282 (c6288_wire_1423, {c6288_wire_1423_0, c6288_wire_1423_1, c6288_wire_1423_2});
fanout_n #(2, 0, 0) FANOUT_283 (c6288_wire_1494, {c6288_wire_1494_0, c6288_wire_1494_1});
fanout_n #(3, 0, 0) FANOUT_284 (c6288_wire_1500, {c6288_wire_1500_0, c6288_wire_1500_1, c6288_wire_1500_2});
fanout_n #(3, 0, 0) FANOUT_285 (c6288_wire_526, {c6288_wire_526_0, c6288_wire_526_1, c6288_wire_526_2});
fanout_n #(2, 0, 0) FANOUT_286 (c6288_wire_1503, {c6288_wire_1503_0, c6288_wire_1503_1});
fanout_n #(3, 0, 0) FANOUT_287 (c6288_wire_524, {c6288_wire_524_0, c6288_wire_524_1, c6288_wire_524_2});
fanout_n #(2, 0, 0) FANOUT_288 (c6288_wire_1509, {c6288_wire_1509_0, c6288_wire_1509_1});
fanout_n #(3, 0, 0) FANOUT_289 (c6288_wire_522, {c6288_wire_522_0, c6288_wire_522_1, c6288_wire_522_2});
fanout_n #(2, 0, 0) FANOUT_290 (c6288_wire_1514, {c6288_wire_1514_0, c6288_wire_1514_1});
fanout_n #(3, 0, 0) FANOUT_291 (c6288_wire_520, {c6288_wire_520_0, c6288_wire_520_1, c6288_wire_520_2});
fanout_n #(2, 0, 0) FANOUT_292 (c6288_wire_1519, {c6288_wire_1519_0, c6288_wire_1519_1});
fanout_n #(3, 0, 0) FANOUT_293 (c6288_wire_518, {c6288_wire_518_0, c6288_wire_518_1, c6288_wire_518_2});
fanout_n #(2, 0, 0) FANOUT_294 (c6288_wire_1524, {c6288_wire_1524_0, c6288_wire_1524_1});
fanout_n #(3, 0, 0) FANOUT_295 (c6288_wire_516, {c6288_wire_516_0, c6288_wire_516_1, c6288_wire_516_2});
fanout_n #(2, 0, 0) FANOUT_296 (c6288_wire_1529, {c6288_wire_1529_0, c6288_wire_1529_1});
fanout_n #(3, 0, 0) FANOUT_297 (c6288_wire_514, {c6288_wire_514_0, c6288_wire_514_1, c6288_wire_514_2});
fanout_n #(2, 0, 0) FANOUT_298 (c6288_wire_1534, {c6288_wire_1534_0, c6288_wire_1534_1});
fanout_n #(3, 0, 0) FANOUT_299 (c6288_wire_512, {c6288_wire_512_0, c6288_wire_512_1, c6288_wire_512_2});
fanout_n #(2, 0, 0) FANOUT_300 (c6288_wire_1539, {c6288_wire_1539_0, c6288_wire_1539_1});
fanout_n #(3, 0, 0) FANOUT_301 (c6288_wire_510, {c6288_wire_510_0, c6288_wire_510_1, c6288_wire_510_2});
fanout_n #(2, 0, 0) FANOUT_302 (c6288_wire_1476, {c6288_wire_1476_0, c6288_wire_1476_1});
fanout_n #(3, 0, 0) FANOUT_303 (c6288_wire_550, {c6288_wire_550_0, c6288_wire_550_1, c6288_wire_550_2});
fanout_n #(2, 0, 0) FANOUT_304 (c6288_wire_1549, {c6288_wire_1549_0, c6288_wire_1549_1});
fanout_n #(3, 0, 0) FANOUT_305 (c6288_wire_548, {c6288_wire_548_0, c6288_wire_548_1, c6288_wire_548_2});
fanout_n #(2, 0, 0) FANOUT_306 (c6288_wire_1557, {c6288_wire_1557_0, c6288_wire_1557_1});
fanout_n #(3, 0, 0) FANOUT_307 (c6288_wire_546, {c6288_wire_546_0, c6288_wire_546_1, c6288_wire_546_2});
fanout_n #(2, 0, 0) FANOUT_308 (c6288_wire_1562, {c6288_wire_1562_0, c6288_wire_1562_1});
fanout_n #(3, 0, 0) FANOUT_309 (c6288_wire_544, {c6288_wire_544_0, c6288_wire_544_1, c6288_wire_544_2});
fanout_n #(2, 0, 0) FANOUT_310 (c6288_wire_1567, {c6288_wire_1567_0, c6288_wire_1567_1});
fanout_n #(3, 0, 0) FANOUT_311 (c6288_wire_1501, {c6288_wire_1501_0, c6288_wire_1501_1, c6288_wire_1501_2});
fanout_n #(2, 0, 0) FANOUT_312 (c6288_wire_1572, {c6288_wire_1572_0, c6288_wire_1572_1});
fanout_n #(3, 0, 0) FANOUT_313 (c6288_wire_1578, {c6288_wire_1578_0, c6288_wire_1578_1, c6288_wire_1578_2});
fanout_n #(3, 0, 0) FANOUT_314 (c6288_wire_568, {c6288_wire_568_0, c6288_wire_568_1, c6288_wire_568_2});
fanout_n #(2, 0, 0) FANOUT_315 (c6288_wire_1581, {c6288_wire_1581_0, c6288_wire_1581_1});
fanout_n #(3, 0, 0) FANOUT_316 (c6288_wire_566, {c6288_wire_566_0, c6288_wire_566_1, c6288_wire_566_2});
fanout_n #(2, 0, 0) FANOUT_317 (c6288_wire_1587, {c6288_wire_1587_0, c6288_wire_1587_1});
fanout_n #(3, 0, 0) FANOUT_318 (c6288_wire_564, {c6288_wire_564_0, c6288_wire_564_1, c6288_wire_564_2});
fanout_n #(2, 0, 0) FANOUT_319 (c6288_wire_1592, {c6288_wire_1592_0, c6288_wire_1592_1});
fanout_n #(3, 0, 0) FANOUT_320 (c6288_wire_562, {c6288_wire_562_0, c6288_wire_562_1, c6288_wire_562_2});
fanout_n #(2, 0, 0) FANOUT_321 (c6288_wire_1597, {c6288_wire_1597_0, c6288_wire_1597_1});
fanout_n #(3, 0, 0) FANOUT_322 (c6288_wire_560, {c6288_wire_560_0, c6288_wire_560_1, c6288_wire_560_2});
fanout_n #(2, 0, 0) FANOUT_323 (c6288_wire_1602, {c6288_wire_1602_0, c6288_wire_1602_1});
fanout_n #(3, 0, 0) FANOUT_324 (c6288_wire_558, {c6288_wire_558_0, c6288_wire_558_1, c6288_wire_558_2});
fanout_n #(2, 0, 0) FANOUT_325 (c6288_wire_1607, {c6288_wire_1607_0, c6288_wire_1607_1});
fanout_n #(3, 0, 0) FANOUT_326 (c6288_wire_556, {c6288_wire_556_0, c6288_wire_556_1, c6288_wire_556_2});
fanout_n #(2, 0, 0) FANOUT_327 (c6288_wire_1612, {c6288_wire_1612_0, c6288_wire_1612_1});
fanout_n #(3, 0, 0) FANOUT_328 (c6288_wire_554, {c6288_wire_554_0, c6288_wire_554_1, c6288_wire_554_2});
fanout_n #(2, 0, 0) FANOUT_329 (c6288_wire_1617, {c6288_wire_1617_0, c6288_wire_1617_1});
fanout_n #(3, 0, 0) FANOUT_330 (c6288_wire_552, {c6288_wire_552_0, c6288_wire_552_1, c6288_wire_552_2});
fanout_n #(2, 0, 0) FANOUT_331 (c6288_wire_1554, {c6288_wire_1554_0, c6288_wire_1554_1});
fanout_n #(3, 0, 0) FANOUT_332 (c6288_wire_592, {c6288_wire_592_0, c6288_wire_592_1, c6288_wire_592_2});
fanout_n #(2, 0, 0) FANOUT_333 (c6288_wire_1627, {c6288_wire_1627_0, c6288_wire_1627_1});
fanout_n #(3, 0, 0) FANOUT_334 (c6288_wire_590, {c6288_wire_590_0, c6288_wire_590_1, c6288_wire_590_2});
fanout_n #(2, 0, 0) FANOUT_335 (c6288_wire_1635, {c6288_wire_1635_0, c6288_wire_1635_1});
fanout_n #(3, 0, 0) FANOUT_336 (c6288_wire_588, {c6288_wire_588_0, c6288_wire_588_1, c6288_wire_588_2});
fanout_n #(2, 0, 0) FANOUT_337 (c6288_wire_1640, {c6288_wire_1640_0, c6288_wire_1640_1});
fanout_n #(3, 0, 0) FANOUT_338 (c6288_wire_586, {c6288_wire_586_0, c6288_wire_586_1, c6288_wire_586_2});
fanout_n #(2, 0, 0) FANOUT_339 (c6288_wire_1645, {c6288_wire_1645_0, c6288_wire_1645_1});
fanout_n #(3, 0, 0) FANOUT_340 (c6288_wire_1579, {c6288_wire_1579_0, c6288_wire_1579_1, c6288_wire_1579_2});
fanout_n #(2, 0, 0) FANOUT_341 (c6288_wire_1650, {c6288_wire_1650_0, c6288_wire_1650_1});
fanout_n #(3, 0, 0) FANOUT_342 (c6288_wire_1656, {c6288_wire_1656_0, c6288_wire_1656_1, c6288_wire_1656_2});
fanout_n #(3, 0, 0) FANOUT_343 (c6288_wire_610, {c6288_wire_610_0, c6288_wire_610_1, c6288_wire_610_2});
fanout_n #(2, 0, 0) FANOUT_344 (c6288_wire_1659, {c6288_wire_1659_0, c6288_wire_1659_1});
fanout_n #(3, 0, 0) FANOUT_345 (c6288_wire_608, {c6288_wire_608_0, c6288_wire_608_1, c6288_wire_608_2});
fanout_n #(2, 0, 0) FANOUT_346 (c6288_wire_1665, {c6288_wire_1665_0, c6288_wire_1665_1});
fanout_n #(3, 0, 0) FANOUT_347 (c6288_wire_606, {c6288_wire_606_0, c6288_wire_606_1, c6288_wire_606_2});
fanout_n #(2, 0, 0) FANOUT_348 (c6288_wire_1670, {c6288_wire_1670_0, c6288_wire_1670_1});
fanout_n #(3, 0, 0) FANOUT_349 (c6288_wire_604, {c6288_wire_604_0, c6288_wire_604_1, c6288_wire_604_2});
fanout_n #(2, 0, 0) FANOUT_350 (c6288_wire_1675, {c6288_wire_1675_0, c6288_wire_1675_1});
fanout_n #(3, 0, 0) FANOUT_351 (c6288_wire_602, {c6288_wire_602_0, c6288_wire_602_1, c6288_wire_602_2});
fanout_n #(2, 0, 0) FANOUT_352 (c6288_wire_1680, {c6288_wire_1680_0, c6288_wire_1680_1});
fanout_n #(3, 0, 0) FANOUT_353 (c6288_wire_600, {c6288_wire_600_0, c6288_wire_600_1, c6288_wire_600_2});
fanout_n #(2, 0, 0) FANOUT_354 (c6288_wire_1685, {c6288_wire_1685_0, c6288_wire_1685_1});
fanout_n #(3, 0, 0) FANOUT_355 (c6288_wire_598, {c6288_wire_598_0, c6288_wire_598_1, c6288_wire_598_2});
fanout_n #(2, 0, 0) FANOUT_356 (c6288_wire_1690, {c6288_wire_1690_0, c6288_wire_1690_1});
fanout_n #(3, 0, 0) FANOUT_357 (c6288_wire_596, {c6288_wire_596_0, c6288_wire_596_1, c6288_wire_596_2});
fanout_n #(2, 0, 0) FANOUT_358 (c6288_wire_1695, {c6288_wire_1695_0, c6288_wire_1695_1});
fanout_n #(3, 0, 0) FANOUT_359 (c6288_wire_594, {c6288_wire_594_0, c6288_wire_594_1, c6288_wire_594_2});
fanout_n #(2, 0, 0) FANOUT_360 (c6288_wire_1632, {c6288_wire_1632_0, c6288_wire_1632_1});
fanout_n #(3, 0, 0) FANOUT_361 (c6288_wire_634, {c6288_wire_634_0, c6288_wire_634_1, c6288_wire_634_2});
fanout_n #(2, 0, 0) FANOUT_362 (c6288_wire_1705, {c6288_wire_1705_0, c6288_wire_1705_1});
fanout_n #(3, 0, 0) FANOUT_363 (c6288_wire_632, {c6288_wire_632_0, c6288_wire_632_1, c6288_wire_632_2});
fanout_n #(2, 0, 0) FANOUT_364 (c6288_wire_1713, {c6288_wire_1713_0, c6288_wire_1713_1});
fanout_n #(3, 0, 0) FANOUT_365 (c6288_wire_630, {c6288_wire_630_0, c6288_wire_630_1, c6288_wire_630_2});
fanout_n #(2, 0, 0) FANOUT_366 (c6288_wire_1718, {c6288_wire_1718_0, c6288_wire_1718_1});
fanout_n #(3, 0, 0) FANOUT_367 (c6288_wire_628, {c6288_wire_628_0, c6288_wire_628_1, c6288_wire_628_2});
fanout_n #(2, 0, 0) FANOUT_368 (c6288_wire_1723, {c6288_wire_1723_0, c6288_wire_1723_1});
fanout_n #(3, 0, 0) FANOUT_369 (c6288_wire_1657, {c6288_wire_1657_0, c6288_wire_1657_1, c6288_wire_1657_2});
fanout_n #(2, 0, 0) FANOUT_370 (c6288_wire_1728, {c6288_wire_1728_0, c6288_wire_1728_1});
fanout_n #(3, 0, 0) FANOUT_371 (c6288_wire_1734, {c6288_wire_1734_0, c6288_wire_1734_1, c6288_wire_1734_2});
fanout_n #(3, 0, 0) FANOUT_372 (c6288_wire_652, {c6288_wire_652_0, c6288_wire_652_1, c6288_wire_652_2});
fanout_n #(2, 0, 0) FANOUT_373 (c6288_wire_1737, {c6288_wire_1737_0, c6288_wire_1737_1});
fanout_n #(3, 0, 0) FANOUT_374 (c6288_wire_650, {c6288_wire_650_0, c6288_wire_650_1, c6288_wire_650_2});
fanout_n #(2, 0, 0) FANOUT_375 (c6288_wire_1743, {c6288_wire_1743_0, c6288_wire_1743_1});
fanout_n #(3, 0, 0) FANOUT_376 (c6288_wire_648, {c6288_wire_648_0, c6288_wire_648_1, c6288_wire_648_2});
fanout_n #(2, 0, 0) FANOUT_377 (c6288_wire_1748, {c6288_wire_1748_0, c6288_wire_1748_1});
fanout_n #(3, 0, 0) FANOUT_378 (c6288_wire_646, {c6288_wire_646_0, c6288_wire_646_1, c6288_wire_646_2});
fanout_n #(2, 0, 0) FANOUT_379 (c6288_wire_1753, {c6288_wire_1753_0, c6288_wire_1753_1});
fanout_n #(3, 0, 0) FANOUT_380 (c6288_wire_644, {c6288_wire_644_0, c6288_wire_644_1, c6288_wire_644_2});
fanout_n #(2, 0, 0) FANOUT_381 (c6288_wire_1758, {c6288_wire_1758_0, c6288_wire_1758_1});
fanout_n #(3, 0, 0) FANOUT_382 (c6288_wire_642, {c6288_wire_642_0, c6288_wire_642_1, c6288_wire_642_2});
fanout_n #(2, 0, 0) FANOUT_383 (c6288_wire_1763, {c6288_wire_1763_0, c6288_wire_1763_1});
fanout_n #(3, 0, 0) FANOUT_384 (c6288_wire_640, {c6288_wire_640_0, c6288_wire_640_1, c6288_wire_640_2});
fanout_n #(2, 0, 0) FANOUT_385 (c6288_wire_1768, {c6288_wire_1768_0, c6288_wire_1768_1});
fanout_n #(3, 0, 0) FANOUT_386 (c6288_wire_638, {c6288_wire_638_0, c6288_wire_638_1, c6288_wire_638_2});
fanout_n #(2, 0, 0) FANOUT_387 (c6288_wire_1773, {c6288_wire_1773_0, c6288_wire_1773_1});
fanout_n #(3, 0, 0) FANOUT_388 (c6288_wire_636, {c6288_wire_636_0, c6288_wire_636_1, c6288_wire_636_2});
fanout_n #(2, 0, 0) FANOUT_389 (c6288_wire_1710, {c6288_wire_1710_0, c6288_wire_1710_1});
fanout_n #(3, 0, 0) FANOUT_390 (c6288_wire_676, {c6288_wire_676_0, c6288_wire_676_1, c6288_wire_676_2});
fanout_n #(2, 0, 0) FANOUT_391 (c6288_wire_1783, {c6288_wire_1783_0, c6288_wire_1783_1});
fanout_n #(3, 0, 0) FANOUT_392 (c6288_wire_674, {c6288_wire_674_0, c6288_wire_674_1, c6288_wire_674_2});
fanout_n #(2, 0, 0) FANOUT_393 (c6288_wire_1791, {c6288_wire_1791_0, c6288_wire_1791_1});
fanout_n #(3, 0, 0) FANOUT_394 (c6288_wire_672, {c6288_wire_672_0, c6288_wire_672_1, c6288_wire_672_2});
fanout_n #(2, 0, 0) FANOUT_395 (c6288_wire_1796, {c6288_wire_1796_0, c6288_wire_1796_1});
fanout_n #(3, 0, 0) FANOUT_396 (c6288_wire_670, {c6288_wire_670_0, c6288_wire_670_1, c6288_wire_670_2});
fanout_n #(2, 0, 0) FANOUT_397 (c6288_wire_1801, {c6288_wire_1801_0, c6288_wire_1801_1});
fanout_n #(3, 0, 0) FANOUT_398 (c6288_wire_1735, {c6288_wire_1735_0, c6288_wire_1735_1, c6288_wire_1735_2});
fanout_n #(2, 0, 0) FANOUT_399 (c6288_wire_1806, {c6288_wire_1806_0, c6288_wire_1806_1});
fanout_n #(3, 0, 0) FANOUT_400 (c6288_wire_1812, {c6288_wire_1812_0, c6288_wire_1812_1, c6288_wire_1812_2});
fanout_n #(3, 0, 0) FANOUT_401 (c6288_wire_694, {c6288_wire_694_0, c6288_wire_694_1, c6288_wire_694_2});
fanout_n #(2, 0, 0) FANOUT_402 (c6288_wire_1815, {c6288_wire_1815_0, c6288_wire_1815_1});
fanout_n #(3, 0, 0) FANOUT_403 (c6288_wire_692, {c6288_wire_692_0, c6288_wire_692_1, c6288_wire_692_2});
fanout_n #(2, 0, 0) FANOUT_404 (c6288_wire_1821, {c6288_wire_1821_0, c6288_wire_1821_1});
fanout_n #(3, 0, 0) FANOUT_405 (c6288_wire_690, {c6288_wire_690_0, c6288_wire_690_1, c6288_wire_690_2});
fanout_n #(2, 0, 0) FANOUT_406 (c6288_wire_1826, {c6288_wire_1826_0, c6288_wire_1826_1});
fanout_n #(3, 0, 0) FANOUT_407 (c6288_wire_688, {c6288_wire_688_0, c6288_wire_688_1, c6288_wire_688_2});
fanout_n #(2, 0, 0) FANOUT_408 (c6288_wire_1831, {c6288_wire_1831_0, c6288_wire_1831_1});
fanout_n #(3, 0, 0) FANOUT_409 (c6288_wire_686, {c6288_wire_686_0, c6288_wire_686_1, c6288_wire_686_2});
fanout_n #(2, 0, 0) FANOUT_410 (c6288_wire_1836, {c6288_wire_1836_0, c6288_wire_1836_1});
fanout_n #(3, 0, 0) FANOUT_411 (c6288_wire_684, {c6288_wire_684_0, c6288_wire_684_1, c6288_wire_684_2});
fanout_n #(2, 0, 0) FANOUT_412 (c6288_wire_1841, {c6288_wire_1841_0, c6288_wire_1841_1});
fanout_n #(3, 0, 0) FANOUT_413 (c6288_wire_682, {c6288_wire_682_0, c6288_wire_682_1, c6288_wire_682_2});
fanout_n #(2, 0, 0) FANOUT_414 (c6288_wire_1846, {c6288_wire_1846_0, c6288_wire_1846_1});
fanout_n #(3, 0, 0) FANOUT_415 (c6288_wire_680, {c6288_wire_680_0, c6288_wire_680_1, c6288_wire_680_2});
fanout_n #(2, 0, 0) FANOUT_416 (c6288_wire_1851, {c6288_wire_1851_0, c6288_wire_1851_1});
fanout_n #(3, 0, 0) FANOUT_417 (c6288_wire_678, {c6288_wire_678_0, c6288_wire_678_1, c6288_wire_678_2});
fanout_n #(2, 0, 0) FANOUT_418 (c6288_wire_1788, {c6288_wire_1788_0, c6288_wire_1788_1});
fanout_n #(3, 0, 0) FANOUT_419 (c6288_wire_718, {c6288_wire_718_0, c6288_wire_718_1, c6288_wire_718_2});
fanout_n #(2, 0, 0) FANOUT_420 (c6288_wire_1861, {c6288_wire_1861_0, c6288_wire_1861_1});
fanout_n #(3, 0, 0) FANOUT_421 (c6288_wire_716, {c6288_wire_716_0, c6288_wire_716_1, c6288_wire_716_2});
fanout_n #(2, 0, 0) FANOUT_422 (c6288_wire_1869, {c6288_wire_1869_0, c6288_wire_1869_1});
fanout_n #(3, 0, 0) FANOUT_423 (c6288_wire_714, {c6288_wire_714_0, c6288_wire_714_1, c6288_wire_714_2});
fanout_n #(2, 0, 0) FANOUT_424 (c6288_wire_1874, {c6288_wire_1874_0, c6288_wire_1874_1});
fanout_n #(3, 0, 0) FANOUT_425 (c6288_wire_712, {c6288_wire_712_0, c6288_wire_712_1, c6288_wire_712_2});
fanout_n #(2, 0, 0) FANOUT_426 (c6288_wire_1879, {c6288_wire_1879_0, c6288_wire_1879_1});
fanout_n #(3, 0, 0) FANOUT_427 (c6288_wire_1813, {c6288_wire_1813_0, c6288_wire_1813_1, c6288_wire_1813_2});
fanout_n #(2, 0, 0) FANOUT_428 (c6288_wire_1884, {c6288_wire_1884_0, c6288_wire_1884_1});
fanout_n #(3, 0, 0) FANOUT_429 (c6288_wire_873, {c6288_wire_873_0, c6288_wire_873_1, c6288_wire_873_2});
fanout_n #(3, 0, 0) FANOUT_430 (c6288_wire_736, {c6288_wire_736_0, c6288_wire_736_1, c6288_wire_736_2});
fanout_n #(2, 0, 0) FANOUT_431 (c6288_wire_1890, {c6288_wire_1890_0, c6288_wire_1890_1});
fanout_n #(3, 0, 0) FANOUT_432 (c6288_wire_734, {c6288_wire_734_0, c6288_wire_734_1, c6288_wire_734_2});
fanout_n #(2, 0, 0) FANOUT_433 (c6288_wire_1896, {c6288_wire_1896_0, c6288_wire_1896_1});
fanout_n #(3, 0, 0) FANOUT_434 (c6288_wire_732, {c6288_wire_732_0, c6288_wire_732_1, c6288_wire_732_2});
fanout_n #(2, 0, 0) FANOUT_435 (c6288_wire_1901, {c6288_wire_1901_0, c6288_wire_1901_1});
fanout_n #(3, 0, 0) FANOUT_436 (c6288_wire_730, {c6288_wire_730_0, c6288_wire_730_1, c6288_wire_730_2});
fanout_n #(2, 0, 0) FANOUT_437 (c6288_wire_1906, {c6288_wire_1906_0, c6288_wire_1906_1});
fanout_n #(3, 0, 0) FANOUT_438 (c6288_wire_728, {c6288_wire_728_0, c6288_wire_728_1, c6288_wire_728_2});
fanout_n #(2, 0, 0) FANOUT_439 (c6288_wire_1911, {c6288_wire_1911_0, c6288_wire_1911_1});
fanout_n #(3, 0, 0) FANOUT_440 (c6288_wire_726, {c6288_wire_726_0, c6288_wire_726_1, c6288_wire_726_2});
fanout_n #(2, 0, 0) FANOUT_441 (c6288_wire_1916, {c6288_wire_1916_0, c6288_wire_1916_1});
fanout_n #(3, 0, 0) FANOUT_442 (c6288_wire_724, {c6288_wire_724_0, c6288_wire_724_1, c6288_wire_724_2});
fanout_n #(2, 0, 0) FANOUT_443 (c6288_wire_1921, {c6288_wire_1921_0, c6288_wire_1921_1});
fanout_n #(3, 0, 0) FANOUT_444 (c6288_wire_722, {c6288_wire_722_0, c6288_wire_722_1, c6288_wire_722_2});
fanout_n #(2, 0, 0) FANOUT_445 (c6288_wire_1926, {c6288_wire_1926_0, c6288_wire_1926_1});
fanout_n #(3, 0, 0) FANOUT_446 (c6288_wire_720, {c6288_wire_720_0, c6288_wire_720_1, c6288_wire_720_2});
fanout_n #(2, 0, 0) FANOUT_447 (c6288_wire_1866, {c6288_wire_1866_0, c6288_wire_1866_1});
fanout_n #(3, 0, 0) FANOUT_448 (c6288_wire_1859, {c6288_wire_1859_0, c6288_wire_1859_1, c6288_wire_1859_2});
fanout_n #(2, 0, 0) FANOUT_449 (c6288_wire_1862, {c6288_wire_1862_0, c6288_wire_1862_1});
fanout_n #(2, 0, 0) FANOUT_450 (c6288_wire_1870, {c6288_wire_1870_0, c6288_wire_1870_1});
fanout_n #(2, 0, 0) FANOUT_451 (c6288_wire_1875, {c6288_wire_1875_0, c6288_wire_1875_1});
fanout_n #(2, 0, 0) FANOUT_452 (c6288_wire_1880, {c6288_wire_1880_0, c6288_wire_1880_1});
fanout_n #(2, 0, 0) FANOUT_453 (c6288_wire_1885, {c6288_wire_1885_0, c6288_wire_1885_1});
fanout_n #(2, 0, 0) FANOUT_454 (c6288_wire_1891, {c6288_wire_1891_0, c6288_wire_1891_1});
fanout_n #(2, 0, 0) FANOUT_455 (c6288_wire_1897, {c6288_wire_1897_0, c6288_wire_1897_1});
fanout_n #(2, 0, 0) FANOUT_456 (c6288_wire_1902, {c6288_wire_1902_0, c6288_wire_1902_1});
fanout_n #(2, 0, 0) FANOUT_457 (c6288_wire_1907, {c6288_wire_1907_0, c6288_wire_1907_1});
fanout_n #(2, 0, 0) FANOUT_458 (c6288_wire_1912, {c6288_wire_1912_0, c6288_wire_1912_1});
fanout_n #(2, 0, 0) FANOUT_459 (c6288_wire_1917, {c6288_wire_1917_0, c6288_wire_1917_1});
fanout_n #(2, 0, 0) FANOUT_460 (c6288_wire_1922, {c6288_wire_1922_0, c6288_wire_1922_1});
fanout_n #(2, 0, 0) FANOUT_461 (c6288_wire_1927, {c6288_wire_1927_0, c6288_wire_1927_1});
fanout_n #(2, 0, 0) FANOUT_462 (c6288_wire_1867, {c6288_wire_1867_0, c6288_wire_1867_1});
fanout_n #(3, 0, 0) FANOUT_463 (c6288_wire_837, {c6288_wire_837_0, c6288_wire_837_1, c6288_wire_837_2});
fanout_n #(2, 0, 0) FANOUT_464 (c6288_wire_840, {c6288_wire_840_0, c6288_wire_840_1});
fanout_n #(2, 0, 0) FANOUT_465 (c6288_wire_848, {c6288_wire_848_0, c6288_wire_848_1});
fanout_n #(2, 0, 0) FANOUT_466 (c6288_wire_853, {c6288_wire_853_0, c6288_wire_853_1});
fanout_n #(2, 0, 0) FANOUT_467 (c6288_wire_858, {c6288_wire_858_0, c6288_wire_858_1});
fanout_n #(2, 0, 0) FANOUT_468 (c6288_wire_864, {c6288_wire_864_0, c6288_wire_864_1});
fanout_n #(2, 0, 0) FANOUT_469 (c6288_wire_875, {c6288_wire_875_0, c6288_wire_875_1});
fanout_n #(2, 0, 0) FANOUT_470 (c6288_wire_881, {c6288_wire_881_0, c6288_wire_881_1});
fanout_n #(2, 0, 0) FANOUT_471 (c6288_wire_886, {c6288_wire_886_0, c6288_wire_886_1});
fanout_n #(2, 0, 0) FANOUT_472 (c6288_wire_891, {c6288_wire_891_0, c6288_wire_891_1});
fanout_n #(2, 0, 0) FANOUT_473 (c6288_wire_896, {c6288_wire_896_0, c6288_wire_896_1});
fanout_n #(2, 0, 0) FANOUT_474 (c6288_wire_901, {c6288_wire_901_0, c6288_wire_901_1});
fanout_n #(2, 0, 0) FANOUT_475 (c6288_wire_906, {c6288_wire_906_0, c6288_wire_906_1});
fanout_n #(2, 0, 0) FANOUT_476 (c6288_wire_911, {c6288_wire_911_0, c6288_wire_911_1});
fanout_n #(2, 0, 0) FANOUT_477 (c6288_wire_845, {c6288_wire_845_0, c6288_wire_845_1});
fanout_n #(3, 0, 0) FANOUT_478 (c6288_wire_918, {c6288_wire_918_0, c6288_wire_918_1, c6288_wire_918_2});
fanout_n #(2, 0, 0) FANOUT_479 (c6288_wire_921, {c6288_wire_921_0, c6288_wire_921_1});
fanout_n #(2, 0, 0) FANOUT_480 (c6288_wire_929, {c6288_wire_929_0, c6288_wire_929_1});
fanout_n #(2, 0, 0) FANOUT_481 (c6288_wire_934, {c6288_wire_934_0, c6288_wire_934_1});
fanout_n #(2, 0, 0) FANOUT_482 (c6288_wire_939, {c6288_wire_939_0, c6288_wire_939_1});
fanout_n #(2, 0, 0) FANOUT_483 (c6288_wire_944, {c6288_wire_944_0, c6288_wire_944_1});
fanout_n #(2, 0, 0) FANOUT_484 (c6288_wire_953, {c6288_wire_953_0, c6288_wire_953_1});
fanout_n #(2, 0, 0) FANOUT_485 (c6288_wire_959, {c6288_wire_959_0, c6288_wire_959_1});
fanout_n #(2, 0, 0) FANOUT_486 (c6288_wire_964, {c6288_wire_964_0, c6288_wire_964_1});
fanout_n #(2, 0, 0) FANOUT_487 (c6288_wire_969, {c6288_wire_969_0, c6288_wire_969_1});
fanout_n #(2, 0, 0) FANOUT_488 (c6288_wire_974, {c6288_wire_974_0, c6288_wire_974_1});
fanout_n #(2, 0, 0) FANOUT_489 (c6288_wire_979, {c6288_wire_979_0, c6288_wire_979_1});
fanout_n #(2, 0, 0) FANOUT_490 (c6288_wire_984, {c6288_wire_984_0, c6288_wire_984_1});
fanout_n #(2, 0, 0) FANOUT_491 (c6288_wire_989, {c6288_wire_989_0, c6288_wire_989_1});
fanout_n #(2, 0, 0) FANOUT_492 (c6288_wire_926, {c6288_wire_926_0, c6288_wire_926_1});
fanout_n #(3, 0, 0) FANOUT_493 (c6288_wire_996, {c6288_wire_996_0, c6288_wire_996_1, c6288_wire_996_2});
fanout_n #(2, 0, 0) FANOUT_494 (c6288_wire_999, {c6288_wire_999_0, c6288_wire_999_1});
fanout_n #(2, 0, 0) FANOUT_495 (c6288_wire_1007, {c6288_wire_1007_0, c6288_wire_1007_1});
fanout_n #(2, 0, 0) FANOUT_496 (c6288_wire_1012, {c6288_wire_1012_0, c6288_wire_1012_1});
fanout_n #(2, 0, 0) FANOUT_497 (c6288_wire_1017, {c6288_wire_1017_0, c6288_wire_1017_1});
fanout_n #(2, 0, 0) FANOUT_498 (c6288_wire_1022, {c6288_wire_1022_0, c6288_wire_1022_1});
fanout_n #(2, 0, 0) FANOUT_499 (c6288_wire_1031, {c6288_wire_1031_0, c6288_wire_1031_1});
fanout_n #(2, 0, 0) FANOUT_500 (c6288_wire_1037, {c6288_wire_1037_0, c6288_wire_1037_1});
fanout_n #(2, 0, 0) FANOUT_501 (c6288_wire_1042, {c6288_wire_1042_0, c6288_wire_1042_1});
fanout_n #(2, 0, 0) FANOUT_502 (c6288_wire_1047, {c6288_wire_1047_0, c6288_wire_1047_1});
fanout_n #(2, 0, 0) FANOUT_503 (c6288_wire_1052, {c6288_wire_1052_0, c6288_wire_1052_1});
fanout_n #(2, 0, 0) FANOUT_504 (c6288_wire_1057, {c6288_wire_1057_0, c6288_wire_1057_1});
fanout_n #(2, 0, 0) FANOUT_505 (c6288_wire_1062, {c6288_wire_1062_0, c6288_wire_1062_1});
fanout_n #(2, 0, 0) FANOUT_506 (c6288_wire_1067, {c6288_wire_1067_0, c6288_wire_1067_1});
fanout_n #(2, 0, 0) FANOUT_507 (c6288_wire_1004, {c6288_wire_1004_0, c6288_wire_1004_1});
fanout_n #(2, 0, 0) FANOUT_508 (c6288_wire_1073, {c6288_wire_1073_0, c6288_wire_1073_1});
fanout_n #(2, 0, 0) FANOUT_509 (c6288_wire_1075, {c6288_wire_1075_0, c6288_wire_1075_1});
fanout_n #(2, 0, 0) FANOUT_510 (c6288_wire_1083, {c6288_wire_1083_0, c6288_wire_1083_1});
fanout_n #(2, 0, 0) FANOUT_511 (c6288_wire_1088, {c6288_wire_1088_0, c6288_wire_1088_1});
fanout_n #(2, 0, 0) FANOUT_512 (c6288_wire_1093, {c6288_wire_1093_0, c6288_wire_1093_1});
fanout_n #(2, 0, 0) FANOUT_513 (c6288_wire_1098, {c6288_wire_1098_0, c6288_wire_1098_1});
fanout_n #(3, 0, 0) FANOUT_514 (c6288_wire_1109, {c6288_wire_1109_0, c6288_wire_1109_1, c6288_wire_1109_2});
fanout_n #(2, 0, 0) FANOUT_515 (c6288_wire_1116, {c6288_wire_1116_0, c6288_wire_1116_1});
fanout_n #(2, 0, 0) FANOUT_516 (c6288_wire_1121, {c6288_wire_1121_0, c6288_wire_1121_1});
fanout_n #(2, 0, 0) FANOUT_517 (c6288_wire_1126, {c6288_wire_1126_0, c6288_wire_1126_1});
fanout_n #(2, 0, 0) FANOUT_518 (c6288_wire_1131, {c6288_wire_1131_0, c6288_wire_1131_1});
fanout_n #(2, 0, 0) FANOUT_519 (c6288_wire_1136, {c6288_wire_1136_0, c6288_wire_1136_1});
fanout_n #(2, 0, 0) FANOUT_520 (c6288_wire_1141, {c6288_wire_1141_0, c6288_wire_1141_1});
fanout_n #(2, 0, 0) FANOUT_521 (c6288_wire_1146, {c6288_wire_1146_0, c6288_wire_1146_1});
fanout_n #(2, 0, 0) FANOUT_522 (c6288_wire_1080, {c6288_wire_1080_0, c6288_wire_1080_1});
fanout_n #(3, 0, 0) FANOUT_523 (c6288_wire_746, {c6288_wire_746_0, c6288_wire_746_1, c6288_wire_746_2});
fanout_n #(2, 0, 0) FANOUT_524 (c6288_wire_750, {c6288_wire_750_0, c6288_wire_750_1});
fanout_n #(2, 0, 0) FANOUT_525 (c6288_wire_759, {c6288_wire_759_0, c6288_wire_759_1});
fanout_n #(2, 0, 0) FANOUT_526 (c6288_wire_765, {c6288_wire_765_0, c6288_wire_765_1});
fanout_n #(2, 0, 0) FANOUT_527 (c6288_wire_771, {c6288_wire_771_0, c6288_wire_771_1});
fanout_n #(2, 0, 0) FANOUT_528 (c6288_wire_777, {c6288_wire_777_0, c6288_wire_777_1});
fanout_n #(2, 0, 0) FANOUT_529 (c6288_wire_786, {c6288_wire_786_0, c6288_wire_786_1});
fanout_n #(2, 0, 0) FANOUT_530 (c6288_wire_793, {c6288_wire_793_0, c6288_wire_793_1});
fanout_n #(2, 0, 0) FANOUT_531 (c6288_wire_799, {c6288_wire_799_0, c6288_wire_799_1});
fanout_n #(2, 0, 0) FANOUT_532 (c6288_wire_805, {c6288_wire_805_0, c6288_wire_805_1});
fanout_n #(2, 0, 0) FANOUT_533 (c6288_wire_811, {c6288_wire_811_0, c6288_wire_811_1});
fanout_n #(2, 0, 0) FANOUT_534 (c6288_wire_817, {c6288_wire_817_0, c6288_wire_817_1});
fanout_n #(2, 0, 0) FANOUT_535 (c6288_wire_823, {c6288_wire_823_0, c6288_wire_823_1});
fanout_n #(2, 0, 0) FANOUT_536 (c6288_wire_829, {c6288_wire_829_0, c6288_wire_829_1});
fanout_n #(2, 0, 0) FANOUT_537 (c6288_wire_755, {c6288_wire_755_0, c6288_wire_755_1});
fanout_n #(3, 0, 0) FANOUT_538 (c6288_wire_1234, {c6288_wire_1234_0, c6288_wire_1234_1, c6288_wire_1234_2});
fanout_n #(2, 0, 0) FANOUT_539 (c6288_wire_1237, {c6288_wire_1237_0, c6288_wire_1237_1});
fanout_n #(2, 0, 0) FANOUT_540 (c6288_wire_1245, {c6288_wire_1245_0, c6288_wire_1245_1});
fanout_n #(2, 0, 0) FANOUT_541 (c6288_wire_1250, {c6288_wire_1250_0, c6288_wire_1250_1});
fanout_n #(2, 0, 0) FANOUT_542 (c6288_wire_1255, {c6288_wire_1255_0, c6288_wire_1255_1});
fanout_n #(2, 0, 0) FANOUT_543 (c6288_wire_1260, {c6288_wire_1260_0, c6288_wire_1260_1});
fanout_n #(2, 0, 0) FANOUT_544 (c6288_wire_1270, {c6288_wire_1270_0, c6288_wire_1270_1});
fanout_n #(2, 0, 0) FANOUT_545 (c6288_wire_1276, {c6288_wire_1276_0, c6288_wire_1276_1});
fanout_n #(2, 0, 0) FANOUT_546 (c6288_wire_1281, {c6288_wire_1281_0, c6288_wire_1281_1});
fanout_n #(2, 0, 0) FANOUT_547 (c6288_wire_1286, {c6288_wire_1286_0, c6288_wire_1286_1});
fanout_n #(2, 0, 0) FANOUT_548 (c6288_wire_1291, {c6288_wire_1291_0, c6288_wire_1291_1});
fanout_n #(2, 0, 0) FANOUT_549 (c6288_wire_1296, {c6288_wire_1296_0, c6288_wire_1296_1});
fanout_n #(2, 0, 0) FANOUT_550 (c6288_wire_1301, {c6288_wire_1301_0, c6288_wire_1301_1});
fanout_n #(2, 0, 0) FANOUT_551 (c6288_wire_1306, {c6288_wire_1306_0, c6288_wire_1306_1});
fanout_n #(2, 0, 0) FANOUT_552 (c6288_wire_1242, {c6288_wire_1242_0, c6288_wire_1242_1});
fanout_n #(3, 0, 0) FANOUT_553 (c6288_wire_1313, {c6288_wire_1313_0, c6288_wire_1313_1, c6288_wire_1313_2});
fanout_n #(2, 0, 0) FANOUT_554 (c6288_wire_1316, {c6288_wire_1316_0, c6288_wire_1316_1});
fanout_n #(2, 0, 0) FANOUT_555 (c6288_wire_1324, {c6288_wire_1324_0, c6288_wire_1324_1});
fanout_n #(2, 0, 0) FANOUT_556 (c6288_wire_1329, {c6288_wire_1329_0, c6288_wire_1329_1});
fanout_n #(2, 0, 0) FANOUT_557 (c6288_wire_1334, {c6288_wire_1334_0, c6288_wire_1334_1});
fanout_n #(2, 0, 0) FANOUT_558 (c6288_wire_1339, {c6288_wire_1339_0, c6288_wire_1339_1});
fanout_n #(2, 0, 0) FANOUT_559 (c6288_wire_1348, {c6288_wire_1348_0, c6288_wire_1348_1});
fanout_n #(2, 0, 0) FANOUT_560 (c6288_wire_1354, {c6288_wire_1354_0, c6288_wire_1354_1});
fanout_n #(2, 0, 0) FANOUT_561 (c6288_wire_1359, {c6288_wire_1359_0, c6288_wire_1359_1});
fanout_n #(2, 0, 0) FANOUT_562 (c6288_wire_1364, {c6288_wire_1364_0, c6288_wire_1364_1});
fanout_n #(2, 0, 0) FANOUT_563 (c6288_wire_1369, {c6288_wire_1369_0, c6288_wire_1369_1});
fanout_n #(2, 0, 0) FANOUT_564 (c6288_wire_1374, {c6288_wire_1374_0, c6288_wire_1374_1});
fanout_n #(2, 0, 0) FANOUT_565 (c6288_wire_1379, {c6288_wire_1379_0, c6288_wire_1379_1});
fanout_n #(2, 0, 0) FANOUT_566 (c6288_wire_1384, {c6288_wire_1384_0, c6288_wire_1384_1});
fanout_n #(2, 0, 0) FANOUT_567 (c6288_wire_1321, {c6288_wire_1321_0, c6288_wire_1321_1});
fanout_n #(3, 0, 0) FANOUT_568 (c6288_wire_1391, {c6288_wire_1391_0, c6288_wire_1391_1, c6288_wire_1391_2});
fanout_n #(2, 0, 0) FANOUT_569 (c6288_wire_1394, {c6288_wire_1394_0, c6288_wire_1394_1});
fanout_n #(2, 0, 0) FANOUT_570 (c6288_wire_1402, {c6288_wire_1402_0, c6288_wire_1402_1});
fanout_n #(2, 0, 0) FANOUT_571 (c6288_wire_1407, {c6288_wire_1407_0, c6288_wire_1407_1});
fanout_n #(2, 0, 0) FANOUT_572 (c6288_wire_1412, {c6288_wire_1412_0, c6288_wire_1412_1});
fanout_n #(2, 0, 0) FANOUT_573 (c6288_wire_1417, {c6288_wire_1417_0, c6288_wire_1417_1});
fanout_n #(2, 0, 0) FANOUT_574 (c6288_wire_1426, {c6288_wire_1426_0, c6288_wire_1426_1});
fanout_n #(2, 0, 0) FANOUT_575 (c6288_wire_1432, {c6288_wire_1432_0, c6288_wire_1432_1});
fanout_n #(2, 0, 0) FANOUT_576 (c6288_wire_1437, {c6288_wire_1437_0, c6288_wire_1437_1});
fanout_n #(2, 0, 0) FANOUT_577 (c6288_wire_1442, {c6288_wire_1442_0, c6288_wire_1442_1});
fanout_n #(2, 0, 0) FANOUT_578 (c6288_wire_1447, {c6288_wire_1447_0, c6288_wire_1447_1});
fanout_n #(2, 0, 0) FANOUT_579 (c6288_wire_1452, {c6288_wire_1452_0, c6288_wire_1452_1});
fanout_n #(2, 0, 0) FANOUT_580 (c6288_wire_1457, {c6288_wire_1457_0, c6288_wire_1457_1});
fanout_n #(2, 0, 0) FANOUT_581 (c6288_wire_1462, {c6288_wire_1462_0, c6288_wire_1462_1});
fanout_n #(2, 0, 0) FANOUT_582 (c6288_wire_1399, {c6288_wire_1399_0, c6288_wire_1399_1});
fanout_n #(3, 0, 0) FANOUT_583 (c6288_wire_1469, {c6288_wire_1469_0, c6288_wire_1469_1, c6288_wire_1469_2});
fanout_n #(2, 0, 0) FANOUT_584 (c6288_wire_1472, {c6288_wire_1472_0, c6288_wire_1472_1});
fanout_n #(2, 0, 0) FANOUT_585 (c6288_wire_1480, {c6288_wire_1480_0, c6288_wire_1480_1});
fanout_n #(2, 0, 0) FANOUT_586 (c6288_wire_1485, {c6288_wire_1485_0, c6288_wire_1485_1});
fanout_n #(2, 0, 0) FANOUT_587 (c6288_wire_1490, {c6288_wire_1490_0, c6288_wire_1490_1});
fanout_n #(2, 0, 0) FANOUT_588 (c6288_wire_1495, {c6288_wire_1495_0, c6288_wire_1495_1});
fanout_n #(2, 0, 0) FANOUT_589 (c6288_wire_1504, {c6288_wire_1504_0, c6288_wire_1504_1});
fanout_n #(2, 0, 0) FANOUT_590 (c6288_wire_1510, {c6288_wire_1510_0, c6288_wire_1510_1});
fanout_n #(2, 0, 0) FANOUT_591 (c6288_wire_1515, {c6288_wire_1515_0, c6288_wire_1515_1});
fanout_n #(2, 0, 0) FANOUT_592 (c6288_wire_1520, {c6288_wire_1520_0, c6288_wire_1520_1});
fanout_n #(2, 0, 0) FANOUT_593 (c6288_wire_1525, {c6288_wire_1525_0, c6288_wire_1525_1});
fanout_n #(2, 0, 0) FANOUT_594 (c6288_wire_1530, {c6288_wire_1530_0, c6288_wire_1530_1});
fanout_n #(2, 0, 0) FANOUT_595 (c6288_wire_1535, {c6288_wire_1535_0, c6288_wire_1535_1});
fanout_n #(2, 0, 0) FANOUT_596 (c6288_wire_1540, {c6288_wire_1540_0, c6288_wire_1540_1});
fanout_n #(2, 0, 0) FANOUT_597 (c6288_wire_1477, {c6288_wire_1477_0, c6288_wire_1477_1});
fanout_n #(3, 0, 0) FANOUT_598 (c6288_wire_1547, {c6288_wire_1547_0, c6288_wire_1547_1, c6288_wire_1547_2});
fanout_n #(2, 0, 0) FANOUT_599 (c6288_wire_1550, {c6288_wire_1550_0, c6288_wire_1550_1});
fanout_n #(2, 0, 0) FANOUT_600 (c6288_wire_1558, {c6288_wire_1558_0, c6288_wire_1558_1});
fanout_n #(2, 0, 0) FANOUT_601 (c6288_wire_1563, {c6288_wire_1563_0, c6288_wire_1563_1});
fanout_n #(2, 0, 0) FANOUT_602 (c6288_wire_1568, {c6288_wire_1568_0, c6288_wire_1568_1});
fanout_n #(2, 0, 0) FANOUT_603 (c6288_wire_1573, {c6288_wire_1573_0, c6288_wire_1573_1});
fanout_n #(2, 0, 0) FANOUT_604 (c6288_wire_1582, {c6288_wire_1582_0, c6288_wire_1582_1});
fanout_n #(2, 0, 0) FANOUT_605 (c6288_wire_1588, {c6288_wire_1588_0, c6288_wire_1588_1});
fanout_n #(2, 0, 0) FANOUT_606 (c6288_wire_1593, {c6288_wire_1593_0, c6288_wire_1593_1});
fanout_n #(2, 0, 0) FANOUT_607 (c6288_wire_1598, {c6288_wire_1598_0, c6288_wire_1598_1});
fanout_n #(2, 0, 0) FANOUT_608 (c6288_wire_1603, {c6288_wire_1603_0, c6288_wire_1603_1});
fanout_n #(2, 0, 0) FANOUT_609 (c6288_wire_1608, {c6288_wire_1608_0, c6288_wire_1608_1});
fanout_n #(2, 0, 0) FANOUT_610 (c6288_wire_1613, {c6288_wire_1613_0, c6288_wire_1613_1});
fanout_n #(2, 0, 0) FANOUT_611 (c6288_wire_1618, {c6288_wire_1618_0, c6288_wire_1618_1});
fanout_n #(2, 0, 0) FANOUT_612 (c6288_wire_1555, {c6288_wire_1555_0, c6288_wire_1555_1});
fanout_n #(3, 0, 0) FANOUT_613 (c6288_wire_1625, {c6288_wire_1625_0, c6288_wire_1625_1, c6288_wire_1625_2});
fanout_n #(2, 0, 0) FANOUT_614 (c6288_wire_1628, {c6288_wire_1628_0, c6288_wire_1628_1});
fanout_n #(2, 0, 0) FANOUT_615 (c6288_wire_1636, {c6288_wire_1636_0, c6288_wire_1636_1});
fanout_n #(2, 0, 0) FANOUT_616 (c6288_wire_1641, {c6288_wire_1641_0, c6288_wire_1641_1});
fanout_n #(2, 0, 0) FANOUT_617 (c6288_wire_1646, {c6288_wire_1646_0, c6288_wire_1646_1});
fanout_n #(2, 0, 0) FANOUT_618 (c6288_wire_1651, {c6288_wire_1651_0, c6288_wire_1651_1});
fanout_n #(2, 0, 0) FANOUT_619 (c6288_wire_1660, {c6288_wire_1660_0, c6288_wire_1660_1});
fanout_n #(2, 0, 0) FANOUT_620 (c6288_wire_1666, {c6288_wire_1666_0, c6288_wire_1666_1});
fanout_n #(2, 0, 0) FANOUT_621 (c6288_wire_1671, {c6288_wire_1671_0, c6288_wire_1671_1});
fanout_n #(2, 0, 0) FANOUT_622 (c6288_wire_1676, {c6288_wire_1676_0, c6288_wire_1676_1});
fanout_n #(2, 0, 0) FANOUT_623 (c6288_wire_1681, {c6288_wire_1681_0, c6288_wire_1681_1});
fanout_n #(2, 0, 0) FANOUT_624 (c6288_wire_1686, {c6288_wire_1686_0, c6288_wire_1686_1});
fanout_n #(2, 0, 0) FANOUT_625 (c6288_wire_1691, {c6288_wire_1691_0, c6288_wire_1691_1});
fanout_n #(2, 0, 0) FANOUT_626 (c6288_wire_1696, {c6288_wire_1696_0, c6288_wire_1696_1});
fanout_n #(2, 0, 0) FANOUT_627 (c6288_wire_1633, {c6288_wire_1633_0, c6288_wire_1633_1});
fanout_n #(3, 0, 0) FANOUT_628 (c6288_wire_1703, {c6288_wire_1703_0, c6288_wire_1703_1, c6288_wire_1703_2});
fanout_n #(2, 0, 0) FANOUT_629 (c6288_wire_1706, {c6288_wire_1706_0, c6288_wire_1706_1});
fanout_n #(2, 0, 0) FANOUT_630 (c6288_wire_1714, {c6288_wire_1714_0, c6288_wire_1714_1});
fanout_n #(2, 0, 0) FANOUT_631 (c6288_wire_1719, {c6288_wire_1719_0, c6288_wire_1719_1});
fanout_n #(2, 0, 0) FANOUT_632 (c6288_wire_1724, {c6288_wire_1724_0, c6288_wire_1724_1});
fanout_n #(2, 0, 0) FANOUT_633 (c6288_wire_1729, {c6288_wire_1729_0, c6288_wire_1729_1});
fanout_n #(2, 0, 0) FANOUT_634 (c6288_wire_1738, {c6288_wire_1738_0, c6288_wire_1738_1});
fanout_n #(2, 0, 0) FANOUT_635 (c6288_wire_1744, {c6288_wire_1744_0, c6288_wire_1744_1});
fanout_n #(2, 0, 0) FANOUT_636 (c6288_wire_1749, {c6288_wire_1749_0, c6288_wire_1749_1});
fanout_n #(2, 0, 0) FANOUT_637 (c6288_wire_1754, {c6288_wire_1754_0, c6288_wire_1754_1});
fanout_n #(2, 0, 0) FANOUT_638 (c6288_wire_1759, {c6288_wire_1759_0, c6288_wire_1759_1});
fanout_n #(2, 0, 0) FANOUT_639 (c6288_wire_1764, {c6288_wire_1764_0, c6288_wire_1764_1});
fanout_n #(2, 0, 0) FANOUT_640 (c6288_wire_1769, {c6288_wire_1769_0, c6288_wire_1769_1});
fanout_n #(2, 0, 0) FANOUT_641 (c6288_wire_1774, {c6288_wire_1774_0, c6288_wire_1774_1});
fanout_n #(2, 0, 0) FANOUT_642 (c6288_wire_1711, {c6288_wire_1711_0, c6288_wire_1711_1});
fanout_n #(3, 0, 0) FANOUT_643 (c6288_wire_1781, {c6288_wire_1781_0, c6288_wire_1781_1, c6288_wire_1781_2});
fanout_n #(2, 0, 0) FANOUT_644 (c6288_wire_1784, {c6288_wire_1784_0, c6288_wire_1784_1});
fanout_n #(2, 0, 0) FANOUT_645 (c6288_wire_1792, {c6288_wire_1792_0, c6288_wire_1792_1});
fanout_n #(2, 0, 0) FANOUT_646 (c6288_wire_1797, {c6288_wire_1797_0, c6288_wire_1797_1});
fanout_n #(2, 0, 0) FANOUT_647 (c6288_wire_1802, {c6288_wire_1802_0, c6288_wire_1802_1});
fanout_n #(2, 0, 0) FANOUT_648 (c6288_wire_1807, {c6288_wire_1807_0, c6288_wire_1807_1});
fanout_n #(2, 0, 0) FANOUT_649 (c6288_wire_1816, {c6288_wire_1816_0, c6288_wire_1816_1});
fanout_n #(2, 0, 0) FANOUT_650 (c6288_wire_1822, {c6288_wire_1822_0, c6288_wire_1822_1});
fanout_n #(2, 0, 0) FANOUT_651 (c6288_wire_1827, {c6288_wire_1827_0, c6288_wire_1827_1});
fanout_n #(2, 0, 0) FANOUT_652 (c6288_wire_1832, {c6288_wire_1832_0, c6288_wire_1832_1});
fanout_n #(2, 0, 0) FANOUT_653 (c6288_wire_1837, {c6288_wire_1837_0, c6288_wire_1837_1});
fanout_n #(2, 0, 0) FANOUT_654 (c6288_wire_1842, {c6288_wire_1842_0, c6288_wire_1842_1});
fanout_n #(2, 0, 0) FANOUT_655 (c6288_wire_1847, {c6288_wire_1847_0, c6288_wire_1847_1});
fanout_n #(2, 0, 0) FANOUT_656 (c6288_wire_1852, {c6288_wire_1852_0, c6288_wire_1852_1});
fanout_n #(2, 0, 0) FANOUT_657 (c6288_wire_1789, {c6288_wire_1789_0, c6288_wire_1789_1});
fanout_n #(3, 0, 0) FANOUT_658 (c6288_wire_2015, {c6288_wire_2015_0, c6288_wire_2015_1, c6288_wire_2015_2});
fanout_n #(3, 0, 0) FANOUT_659 (c6288_wire_160, {c6288_wire_160_0, c6288_wire_160_1, c6288_wire_160_2});
fanout_n #(3, 0, 0) FANOUT_660 (c6288_wire_202, {c6288_wire_202_0, c6288_wire_202_1, c6288_wire_202_2});
fanout_n #(3, 0, 0) FANOUT_661 (c6288_wire_244, {c6288_wire_244_0, c6288_wire_244_1, c6288_wire_244_2});
fanout_n #(3, 0, 0) FANOUT_662 (c6288_wire_284, {c6288_wire_284_0, c6288_wire_284_1, c6288_wire_284_2});
fanout_n #(3, 0, 0) FANOUT_663 (c6288_wire_311, {c6288_wire_311_0, c6288_wire_311_1, c6288_wire_311_2});
fanout_n #(3, 0, 0) FANOUT_664 (c6288_wire_309, {c6288_wire_309_0, c6288_wire_309_1, c6288_wire_309_2});
fanout_n #(3, 0, 0) FANOUT_665 (c6288_wire_307, {c6288_wire_307_0, c6288_wire_307_1, c6288_wire_307_2});
fanout_n #(3, 0, 0) FANOUT_666 (c6288_wire_305, {c6288_wire_305_0, c6288_wire_305_1, c6288_wire_305_2});
fanout_n #(3, 0, 0) FANOUT_667 (c6288_wire_303, {c6288_wire_303_0, c6288_wire_303_1, c6288_wire_303_2});
fanout_n #(2, 0, 0) FANOUT_668 (c6288_wire_1104, {c6288_wire_1104_0, c6288_wire_1104_1});
fanout_n #(3, 0, 0) FANOUT_669 (c6288_wire_2230, {c6288_wire_2230_0, c6288_wire_2230_1, c6288_wire_2230_2});
fanout_n #(3, 0, 0) FANOUT_670 (c6288_wire_325, {c6288_wire_325_0, c6288_wire_325_1, c6288_wire_325_2});
fanout_n #(3, 0, 0) FANOUT_671 (c6288_wire_323, {c6288_wire_323_0, c6288_wire_323_1, c6288_wire_323_2});
fanout_n #(3, 0, 0) FANOUT_672 (c6288_wire_321, {c6288_wire_321_0, c6288_wire_321_1, c6288_wire_321_2});
fanout_n #(3, 0, 0) FANOUT_673 (c6288_wire_319, {c6288_wire_319_0, c6288_wire_319_1, c6288_wire_319_2});
fanout_n #(3, 0, 0) FANOUT_674 (c6288_wire_317, {c6288_wire_317_0, c6288_wire_317_1, c6288_wire_317_2});
fanout_n #(3, 0, 0) FANOUT_675 (c6288_wire_315, {c6288_wire_315_0, c6288_wire_315_1, c6288_wire_315_2});
fanout_n #(3, 0, 0) FANOUT_676 (c6288_wire_313, {c6288_wire_313_0, c6288_wire_313_1, c6288_wire_313_2});
fanout_n #(3, 0, 0) FANOUT_677 (c6288_wire_402, {c6288_wire_402_0, c6288_wire_402_1, c6288_wire_402_2});
fanout_n #(3, 0, 0) FANOUT_678 (c6288_wire_444, {c6288_wire_444_0, c6288_wire_444_1, c6288_wire_444_2});
fanout_n #(3, 0, 0) FANOUT_679 (c6288_wire_486, {c6288_wire_486_0, c6288_wire_486_1, c6288_wire_486_2});
fanout_n #(3, 0, 0) FANOUT_680 (c6288_wire_528, {c6288_wire_528_0, c6288_wire_528_1, c6288_wire_528_2});
fanout_n #(3, 0, 0) FANOUT_681 (c6288_wire_570, {c6288_wire_570_0, c6288_wire_570_1, c6288_wire_570_2});
fanout_n #(3, 0, 0) FANOUT_682 (c6288_wire_612, {c6288_wire_612_0, c6288_wire_612_1, c6288_wire_612_2});
fanout_n #(3, 0, 0) FANOUT_683 (c6288_wire_654, {c6288_wire_654_0, c6288_wire_654_1, c6288_wire_654_2});
fanout_n #(3, 0, 0) FANOUT_684 (c6288_wire_696, {c6288_wire_696_0, c6288_wire_696_1, c6288_wire_696_2});
fanout_n #(3, 0, 0) FANOUT_685 (c6288_wire_738, {c6288_wire_738_0, c6288_wire_738_1, c6288_wire_738_2});
fanout_n #(2, 0, 0) FANOUT_686 (c6288_wire_756, {c6288_wire_756_0, c6288_wire_756_1});
fanout_n #(2, 0, 0) FANOUT_687 (c6288_wire_762, {c6288_wire_762_0, c6288_wire_762_1});
fanout_n #(2, 0, 0) FANOUT_688 (c6288_wire_768, {c6288_wire_768_0, c6288_wire_768_1});
fanout_n #(2, 0, 0) FANOUT_689 (c6288_wire_774, {c6288_wire_774_0, c6288_wire_774_1});
fanout_n #(2, 0, 0) FANOUT_690 (c6288_wire_779, {c6288_wire_779_0, c6288_wire_779_1});
fanout_n #(2, 0, 0) FANOUT_691 (c6288_wire_790, {c6288_wire_790_0, c6288_wire_790_1});
fanout_n #(2, 0, 0) FANOUT_692 (c6288_wire_796, {c6288_wire_796_0, c6288_wire_796_1});
fanout_n #(2, 0, 0) FANOUT_693 (c6288_wire_802, {c6288_wire_802_0, c6288_wire_802_1});
fanout_n #(2, 0, 0) FANOUT_694 (c6288_wire_808, {c6288_wire_808_0, c6288_wire_808_1});
fanout_n #(2, 0, 0) FANOUT_695 (c6288_wire_814, {c6288_wire_814_0, c6288_wire_814_1});
fanout_n #(2, 0, 0) FANOUT_696 (c6288_wire_820, {c6288_wire_820_0, c6288_wire_820_1});
fanout_n #(2, 0, 0) FANOUT_697 (c6288_wire_826, {c6288_wire_826_0, c6288_wire_826_1});
fanout_n #(2, 0, 0) FANOUT_698 (c6288_wire_832, {c6288_wire_832_0, c6288_wire_832_1});
fanout_n #(2, 0, 0) FANOUT_699 (c6288_wire_835, {c6288_wire_835_0, c6288_wire_835_1});
fanout_n #(4, 0, 0) FANOUT_700 (c6288_wire_740, {c6288_wire_740_0, c6288_wire_740_1, c6288_wire_740_2, c6288_wire_740_3});
fanout_n #(32, 0, 0) FANOUT_701 (c6288_wire_32, {c6288_wire_32_0, c6288_wire_32_1, c6288_wire_32_2, c6288_wire_32_3, c6288_wire_32_4, c6288_wire_32_5, c6288_wire_32_6, c6288_wire_32_7, c6288_wire_32_8, c6288_wire_32_9, c6288_wire_32_10, c6288_wire_32_11, c6288_wire_32_12, c6288_wire_32_13, c6288_wire_32_14, c6288_wire_32_15, c6288_wire_32_16, c6288_wire_32_17, c6288_wire_32_18, c6288_wire_32_19, c6288_wire_32_20, c6288_wire_32_21, c6288_wire_32_22, c6288_wire_32_23, c6288_wire_32_24, c6288_wire_32_25, c6288_wire_32_26, c6288_wire_32_27, c6288_wire_32_28, c6288_wire_32_29, c6288_wire_32_30, c6288_wire_32_31});
fanout_n #(46, 0, 0) FANOUT_702 (c6288_wire_57, {c6288_wire_57_0, c6288_wire_57_1, c6288_wire_57_2, c6288_wire_57_3, c6288_wire_57_4, c6288_wire_57_5, c6288_wire_57_6, c6288_wire_57_7, c6288_wire_57_8, c6288_wire_57_9, c6288_wire_57_10, c6288_wire_57_11, c6288_wire_57_12, c6288_wire_57_13, c6288_wire_57_14, c6288_wire_57_15, c6288_wire_57_16, c6288_wire_57_17, c6288_wire_57_18, c6288_wire_57_19, c6288_wire_57_20, c6288_wire_57_21, c6288_wire_57_22, c6288_wire_57_23, c6288_wire_57_24, c6288_wire_57_25, c6288_wire_57_26, c6288_wire_57_27, c6288_wire_57_28, c6288_wire_57_29, c6288_wire_57_30, c6288_wire_57_31, c6288_wire_57_32, c6288_wire_57_33, c6288_wire_57_34, c6288_wire_57_35, c6288_wire_57_36, c6288_wire_57_37, c6288_wire_57_38, c6288_wire_57_39, c6288_wire_57_40, c6288_wire_57_41, c6288_wire_57_42, c6288_wire_57_43, c6288_wire_57_44, c6288_wire_57_45});
fanout_n #(46, 0, 0) FANOUT_703 (c6288_wire_62, {c6288_wire_62_0, c6288_wire_62_1, c6288_wire_62_2, c6288_wire_62_3, c6288_wire_62_4, c6288_wire_62_5, c6288_wire_62_6, c6288_wire_62_7, c6288_wire_62_8, c6288_wire_62_9, c6288_wire_62_10, c6288_wire_62_11, c6288_wire_62_12, c6288_wire_62_13, c6288_wire_62_14, c6288_wire_62_15, c6288_wire_62_16, c6288_wire_62_17, c6288_wire_62_18, c6288_wire_62_19, c6288_wire_62_20, c6288_wire_62_21, c6288_wire_62_22, c6288_wire_62_23, c6288_wire_62_24, c6288_wire_62_25, c6288_wire_62_26, c6288_wire_62_27, c6288_wire_62_28, c6288_wire_62_29, c6288_wire_62_30, c6288_wire_62_31, c6288_wire_62_32, c6288_wire_62_33, c6288_wire_62_34, c6288_wire_62_35, c6288_wire_62_36, c6288_wire_62_37, c6288_wire_62_38, c6288_wire_62_39, c6288_wire_62_40, c6288_wire_62_41, c6288_wire_62_42, c6288_wire_62_43, c6288_wire_62_44, c6288_wire_62_45});
fanout_n #(46, 0, 0) FANOUT_704 (c6288_wire_67, {c6288_wire_67_0, c6288_wire_67_1, c6288_wire_67_2, c6288_wire_67_3, c6288_wire_67_4, c6288_wire_67_5, c6288_wire_67_6, c6288_wire_67_7, c6288_wire_67_8, c6288_wire_67_9, c6288_wire_67_10, c6288_wire_67_11, c6288_wire_67_12, c6288_wire_67_13, c6288_wire_67_14, c6288_wire_67_15, c6288_wire_67_16, c6288_wire_67_17, c6288_wire_67_18, c6288_wire_67_19, c6288_wire_67_20, c6288_wire_67_21, c6288_wire_67_22, c6288_wire_67_23, c6288_wire_67_24, c6288_wire_67_25, c6288_wire_67_26, c6288_wire_67_27, c6288_wire_67_28, c6288_wire_67_29, c6288_wire_67_30, c6288_wire_67_31, c6288_wire_67_32, c6288_wire_67_33, c6288_wire_67_34, c6288_wire_67_35, c6288_wire_67_36, c6288_wire_67_37, c6288_wire_67_38, c6288_wire_67_39, c6288_wire_67_40, c6288_wire_67_41, c6288_wire_67_42, c6288_wire_67_43, c6288_wire_67_44, c6288_wire_67_45});
fanout_n #(46, 0, 0) FANOUT_705 (c6288_wire_5, {c6288_wire_5_0, c6288_wire_5_1, c6288_wire_5_2, c6288_wire_5_3, c6288_wire_5_4, c6288_wire_5_5, c6288_wire_5_6, c6288_wire_5_7, c6288_wire_5_8, c6288_wire_5_9, c6288_wire_5_10, c6288_wire_5_11, c6288_wire_5_12, c6288_wire_5_13, c6288_wire_5_14, c6288_wire_5_15, c6288_wire_5_16, c6288_wire_5_17, c6288_wire_5_18, c6288_wire_5_19, c6288_wire_5_20, c6288_wire_5_21, c6288_wire_5_22, c6288_wire_5_23, c6288_wire_5_24, c6288_wire_5_25, c6288_wire_5_26, c6288_wire_5_27, c6288_wire_5_28, c6288_wire_5_29, c6288_wire_5_30, c6288_wire_5_31, c6288_wire_5_32, c6288_wire_5_33, c6288_wire_5_34, c6288_wire_5_35, c6288_wire_5_36, c6288_wire_5_37, c6288_wire_5_38, c6288_wire_5_39, c6288_wire_5_40, c6288_wire_5_41, c6288_wire_5_42, c6288_wire_5_43, c6288_wire_5_44, c6288_wire_5_45});
fanout_n #(46, 0, 0) FANOUT_706 (c6288_wire_2, {c6288_wire_2_0, c6288_wire_2_1, c6288_wire_2_2, c6288_wire_2_3, c6288_wire_2_4, c6288_wire_2_5, c6288_wire_2_6, c6288_wire_2_7, c6288_wire_2_8, c6288_wire_2_9, c6288_wire_2_10, c6288_wire_2_11, c6288_wire_2_12, c6288_wire_2_13, c6288_wire_2_14, c6288_wire_2_15, c6288_wire_2_16, c6288_wire_2_17, c6288_wire_2_18, c6288_wire_2_19, c6288_wire_2_20, c6288_wire_2_21, c6288_wire_2_22, c6288_wire_2_23, c6288_wire_2_24, c6288_wire_2_25, c6288_wire_2_26, c6288_wire_2_27, c6288_wire_2_28, c6288_wire_2_29, c6288_wire_2_30, c6288_wire_2_31, c6288_wire_2_32, c6288_wire_2_33, c6288_wire_2_34, c6288_wire_2_35, c6288_wire_2_36, c6288_wire_2_37, c6288_wire_2_38, c6288_wire_2_39, c6288_wire_2_40, c6288_wire_2_41, c6288_wire_2_42, c6288_wire_2_43, c6288_wire_2_44, c6288_wire_2_45});
fanout_n #(46, 0, 0) FANOUT_707 (c6288_wire_30, {c6288_wire_30_0, c6288_wire_30_1, c6288_wire_30_2, c6288_wire_30_3, c6288_wire_30_4, c6288_wire_30_5, c6288_wire_30_6, c6288_wire_30_7, c6288_wire_30_8, c6288_wire_30_9, c6288_wire_30_10, c6288_wire_30_11, c6288_wire_30_12, c6288_wire_30_13, c6288_wire_30_14, c6288_wire_30_15, c6288_wire_30_16, c6288_wire_30_17, c6288_wire_30_18, c6288_wire_30_19, c6288_wire_30_20, c6288_wire_30_21, c6288_wire_30_22, c6288_wire_30_23, c6288_wire_30_24, c6288_wire_30_25, c6288_wire_30_26, c6288_wire_30_27, c6288_wire_30_28, c6288_wire_30_29, c6288_wire_30_30, c6288_wire_30_31, c6288_wire_30_32, c6288_wire_30_33, c6288_wire_30_34, c6288_wire_30_35, c6288_wire_30_36, c6288_wire_30_37, c6288_wire_30_38, c6288_wire_30_39, c6288_wire_30_40, c6288_wire_30_41, c6288_wire_30_42, c6288_wire_30_43, c6288_wire_30_44, c6288_wire_30_45});
fanout_n #(46, 0, 0) FANOUT_708 (c6288_wire_10, {c6288_wire_10_0, c6288_wire_10_1, c6288_wire_10_2, c6288_wire_10_3, c6288_wire_10_4, c6288_wire_10_5, c6288_wire_10_6, c6288_wire_10_7, c6288_wire_10_8, c6288_wire_10_9, c6288_wire_10_10, c6288_wire_10_11, c6288_wire_10_12, c6288_wire_10_13, c6288_wire_10_14, c6288_wire_10_15, c6288_wire_10_16, c6288_wire_10_17, c6288_wire_10_18, c6288_wire_10_19, c6288_wire_10_20, c6288_wire_10_21, c6288_wire_10_22, c6288_wire_10_23, c6288_wire_10_24, c6288_wire_10_25, c6288_wire_10_26, c6288_wire_10_27, c6288_wire_10_28, c6288_wire_10_29, c6288_wire_10_30, c6288_wire_10_31, c6288_wire_10_32, c6288_wire_10_33, c6288_wire_10_34, c6288_wire_10_35, c6288_wire_10_36, c6288_wire_10_37, c6288_wire_10_38, c6288_wire_10_39, c6288_wire_10_40, c6288_wire_10_41, c6288_wire_10_42, c6288_wire_10_43, c6288_wire_10_44, c6288_wire_10_45});
fanout_n #(46, 0, 0) FANOUT_709 (c6288_wire_15, {c6288_wire_15_0, c6288_wire_15_1, c6288_wire_15_2, c6288_wire_15_3, c6288_wire_15_4, c6288_wire_15_5, c6288_wire_15_6, c6288_wire_15_7, c6288_wire_15_8, c6288_wire_15_9, c6288_wire_15_10, c6288_wire_15_11, c6288_wire_15_12, c6288_wire_15_13, c6288_wire_15_14, c6288_wire_15_15, c6288_wire_15_16, c6288_wire_15_17, c6288_wire_15_18, c6288_wire_15_19, c6288_wire_15_20, c6288_wire_15_21, c6288_wire_15_22, c6288_wire_15_23, c6288_wire_15_24, c6288_wire_15_25, c6288_wire_15_26, c6288_wire_15_27, c6288_wire_15_28, c6288_wire_15_29, c6288_wire_15_30, c6288_wire_15_31, c6288_wire_15_32, c6288_wire_15_33, c6288_wire_15_34, c6288_wire_15_35, c6288_wire_15_36, c6288_wire_15_37, c6288_wire_15_38, c6288_wire_15_39, c6288_wire_15_40, c6288_wire_15_41, c6288_wire_15_42, c6288_wire_15_43, c6288_wire_15_44, c6288_wire_15_45});
fanout_n #(46, 0, 0) FANOUT_710 (c6288_wire_20, {c6288_wire_20_0, c6288_wire_20_1, c6288_wire_20_2, c6288_wire_20_3, c6288_wire_20_4, c6288_wire_20_5, c6288_wire_20_6, c6288_wire_20_7, c6288_wire_20_8, c6288_wire_20_9, c6288_wire_20_10, c6288_wire_20_11, c6288_wire_20_12, c6288_wire_20_13, c6288_wire_20_14, c6288_wire_20_15, c6288_wire_20_16, c6288_wire_20_17, c6288_wire_20_18, c6288_wire_20_19, c6288_wire_20_20, c6288_wire_20_21, c6288_wire_20_22, c6288_wire_20_23, c6288_wire_20_24, c6288_wire_20_25, c6288_wire_20_26, c6288_wire_20_27, c6288_wire_20_28, c6288_wire_20_29, c6288_wire_20_30, c6288_wire_20_31, c6288_wire_20_32, c6288_wire_20_33, c6288_wire_20_34, c6288_wire_20_35, c6288_wire_20_36, c6288_wire_20_37, c6288_wire_20_38, c6288_wire_20_39, c6288_wire_20_40, c6288_wire_20_41, c6288_wire_20_42, c6288_wire_20_43, c6288_wire_20_44, c6288_wire_20_45});
fanout_n #(45, 0, 0) FANOUT_711 (c6288_wire_25, {c6288_wire_25_0, c6288_wire_25_1, c6288_wire_25_2, c6288_wire_25_3, c6288_wire_25_4, c6288_wire_25_5, c6288_wire_25_6, c6288_wire_25_7, c6288_wire_25_8, c6288_wire_25_9, c6288_wire_25_10, c6288_wire_25_11, c6288_wire_25_12, c6288_wire_25_13, c6288_wire_25_14, c6288_wire_25_15, c6288_wire_25_16, c6288_wire_25_17, c6288_wire_25_18, c6288_wire_25_19, c6288_wire_25_20, c6288_wire_25_21, c6288_wire_25_22, c6288_wire_25_23, c6288_wire_25_24, c6288_wire_25_25, c6288_wire_25_26, c6288_wire_25_27, c6288_wire_25_28, c6288_wire_25_29, c6288_wire_25_30, c6288_wire_25_31, c6288_wire_25_32, c6288_wire_25_33, c6288_wire_25_34, c6288_wire_25_35, c6288_wire_25_36, c6288_wire_25_37, c6288_wire_25_38, c6288_wire_25_39, c6288_wire_25_40, c6288_wire_25_41, c6288_wire_25_42, c6288_wire_25_43, c6288_wire_25_44});
fanout_n #(44, 0, 0) FANOUT_712 (c6288_wire_330, {c6288_wire_330_0, c6288_wire_330_1, c6288_wire_330_2, c6288_wire_330_3, c6288_wire_330_4, c6288_wire_330_5, c6288_wire_330_6, c6288_wire_330_7, c6288_wire_330_8, c6288_wire_330_9, c6288_wire_330_10, c6288_wire_330_11, c6288_wire_330_12, c6288_wire_330_13, c6288_wire_330_14, c6288_wire_330_15, c6288_wire_330_16, c6288_wire_330_17, c6288_wire_330_18, c6288_wire_330_19, c6288_wire_330_20, c6288_wire_330_21, c6288_wire_330_22, c6288_wire_330_23, c6288_wire_330_24, c6288_wire_330_25, c6288_wire_330_26, c6288_wire_330_27, c6288_wire_330_28, c6288_wire_330_29, c6288_wire_330_30, c6288_wire_330_31, c6288_wire_330_32, c6288_wire_330_33, c6288_wire_330_34, c6288_wire_330_35, c6288_wire_330_36, c6288_wire_330_37, c6288_wire_330_38, c6288_wire_330_39, c6288_wire_330_40, c6288_wire_330_41, c6288_wire_330_42, c6288_wire_330_43});
fanout_n #(18, 0, 0) FANOUT_713 (c6288_wire_3, {c6288_wire_3_0, c6288_wire_3_1, c6288_wire_3_2, c6288_wire_3_3, c6288_wire_3_4, c6288_wire_3_5, c6288_wire_3_6, c6288_wire_3_7, c6288_wire_3_8, c6288_wire_3_9, c6288_wire_3_10, c6288_wire_3_11, c6288_wire_3_12, c6288_wire_3_13, c6288_wire_3_14, c6288_wire_3_15, c6288_wire_3_16, c6288_wire_3_17});
fanout_n #(48, 0, 0) FANOUT_714 (c6288_wire_6, {c6288_wire_6_0, c6288_wire_6_1, c6288_wire_6_2, c6288_wire_6_3, c6288_wire_6_4, c6288_wire_6_5, c6288_wire_6_6, c6288_wire_6_7, c6288_wire_6_8, c6288_wire_6_9, c6288_wire_6_10, c6288_wire_6_11, c6288_wire_6_12, c6288_wire_6_13, c6288_wire_6_14, c6288_wire_6_15, c6288_wire_6_16, c6288_wire_6_17, c6288_wire_6_18, c6288_wire_6_19, c6288_wire_6_20, c6288_wire_6_21, c6288_wire_6_22, c6288_wire_6_23, c6288_wire_6_24, c6288_wire_6_25, c6288_wire_6_26, c6288_wire_6_27, c6288_wire_6_28, c6288_wire_6_29, c6288_wire_6_30, c6288_wire_6_31, c6288_wire_6_32, c6288_wire_6_33, c6288_wire_6_34, c6288_wire_6_35, c6288_wire_6_36, c6288_wire_6_37, c6288_wire_6_38, c6288_wire_6_39, c6288_wire_6_40, c6288_wire_6_41, c6288_wire_6_42, c6288_wire_6_43, c6288_wire_6_44, c6288_wire_6_45, c6288_wire_6_46, c6288_wire_6_47});
fanout_n #(46, 0, 0) FANOUT_715 (c6288_wire_78, {c6288_wire_78_0, c6288_wire_78_1, c6288_wire_78_2, c6288_wire_78_3, c6288_wire_78_4, c6288_wire_78_5, c6288_wire_78_6, c6288_wire_78_7, c6288_wire_78_8, c6288_wire_78_9, c6288_wire_78_10, c6288_wire_78_11, c6288_wire_78_12, c6288_wire_78_13, c6288_wire_78_14, c6288_wire_78_15, c6288_wire_78_16, c6288_wire_78_17, c6288_wire_78_18, c6288_wire_78_19, c6288_wire_78_20, c6288_wire_78_21, c6288_wire_78_22, c6288_wire_78_23, c6288_wire_78_24, c6288_wire_78_25, c6288_wire_78_26, c6288_wire_78_27, c6288_wire_78_28, c6288_wire_78_29, c6288_wire_78_30, c6288_wire_78_31, c6288_wire_78_32, c6288_wire_78_33, c6288_wire_78_34, c6288_wire_78_35, c6288_wire_78_36, c6288_wire_78_37, c6288_wire_78_38, c6288_wire_78_39, c6288_wire_78_40, c6288_wire_78_41, c6288_wire_78_42, c6288_wire_78_43, c6288_wire_78_44, c6288_wire_78_45});
fanout_n #(47, 0, 0) FANOUT_716 (c6288_wire_81, {c6288_wire_81_0, c6288_wire_81_1, c6288_wire_81_2, c6288_wire_81_3, c6288_wire_81_4, c6288_wire_81_5, c6288_wire_81_6, c6288_wire_81_7, c6288_wire_81_8, c6288_wire_81_9, c6288_wire_81_10, c6288_wire_81_11, c6288_wire_81_12, c6288_wire_81_13, c6288_wire_81_14, c6288_wire_81_15, c6288_wire_81_16, c6288_wire_81_17, c6288_wire_81_18, c6288_wire_81_19, c6288_wire_81_20, c6288_wire_81_21, c6288_wire_81_22, c6288_wire_81_23, c6288_wire_81_24, c6288_wire_81_25, c6288_wire_81_26, c6288_wire_81_27, c6288_wire_81_28, c6288_wire_81_29, c6288_wire_81_30, c6288_wire_81_31, c6288_wire_81_32, c6288_wire_81_33, c6288_wire_81_34, c6288_wire_81_35, c6288_wire_81_36, c6288_wire_81_37, c6288_wire_81_38, c6288_wire_81_39, c6288_wire_81_40, c6288_wire_81_41, c6288_wire_81_42, c6288_wire_81_43, c6288_wire_81_44, c6288_wire_81_45, c6288_wire_81_46});
fanout_n #(47, 0, 0) FANOUT_717 (c6288_wire_84, {c6288_wire_84_0, c6288_wire_84_1, c6288_wire_84_2, c6288_wire_84_3, c6288_wire_84_4, c6288_wire_84_5, c6288_wire_84_6, c6288_wire_84_7, c6288_wire_84_8, c6288_wire_84_9, c6288_wire_84_10, c6288_wire_84_11, c6288_wire_84_12, c6288_wire_84_13, c6288_wire_84_14, c6288_wire_84_15, c6288_wire_84_16, c6288_wire_84_17, c6288_wire_84_18, c6288_wire_84_19, c6288_wire_84_20, c6288_wire_84_21, c6288_wire_84_22, c6288_wire_84_23, c6288_wire_84_24, c6288_wire_84_25, c6288_wire_84_26, c6288_wire_84_27, c6288_wire_84_28, c6288_wire_84_29, c6288_wire_84_30, c6288_wire_84_31, c6288_wire_84_32, c6288_wire_84_33, c6288_wire_84_34, c6288_wire_84_35, c6288_wire_84_36, c6288_wire_84_37, c6288_wire_84_38, c6288_wire_84_39, c6288_wire_84_40, c6288_wire_84_41, c6288_wire_84_42, c6288_wire_84_43, c6288_wire_84_44, c6288_wire_84_45, c6288_wire_84_46});
fanout_n #(46, 0, 0) FANOUT_718 (c6288_wire_37, {c6288_wire_37_0, c6288_wire_37_1, c6288_wire_37_2, c6288_wire_37_3, c6288_wire_37_4, c6288_wire_37_5, c6288_wire_37_6, c6288_wire_37_7, c6288_wire_37_8, c6288_wire_37_9, c6288_wire_37_10, c6288_wire_37_11, c6288_wire_37_12, c6288_wire_37_13, c6288_wire_37_14, c6288_wire_37_15, c6288_wire_37_16, c6288_wire_37_17, c6288_wire_37_18, c6288_wire_37_19, c6288_wire_37_20, c6288_wire_37_21, c6288_wire_37_22, c6288_wire_37_23, c6288_wire_37_24, c6288_wire_37_25, c6288_wire_37_26, c6288_wire_37_27, c6288_wire_37_28, c6288_wire_37_29, c6288_wire_37_30, c6288_wire_37_31, c6288_wire_37_32, c6288_wire_37_33, c6288_wire_37_34, c6288_wire_37_35, c6288_wire_37_36, c6288_wire_37_37, c6288_wire_37_38, c6288_wire_37_39, c6288_wire_37_40, c6288_wire_37_41, c6288_wire_37_42, c6288_wire_37_43, c6288_wire_37_44, c6288_wire_37_45});
fanout_n #(47, 0, 0) FANOUT_719 (c6288_wire_87, {c6288_wire_87_0, c6288_wire_87_1, c6288_wire_87_2, c6288_wire_87_3, c6288_wire_87_4, c6288_wire_87_5, c6288_wire_87_6, c6288_wire_87_7, c6288_wire_87_8, c6288_wire_87_9, c6288_wire_87_10, c6288_wire_87_11, c6288_wire_87_12, c6288_wire_87_13, c6288_wire_87_14, c6288_wire_87_15, c6288_wire_87_16, c6288_wire_87_17, c6288_wire_87_18, c6288_wire_87_19, c6288_wire_87_20, c6288_wire_87_21, c6288_wire_87_22, c6288_wire_87_23, c6288_wire_87_24, c6288_wire_87_25, c6288_wire_87_26, c6288_wire_87_27, c6288_wire_87_28, c6288_wire_87_29, c6288_wire_87_30, c6288_wire_87_31, c6288_wire_87_32, c6288_wire_87_33, c6288_wire_87_34, c6288_wire_87_35, c6288_wire_87_36, c6288_wire_87_37, c6288_wire_87_38, c6288_wire_87_39, c6288_wire_87_40, c6288_wire_87_41, c6288_wire_87_42, c6288_wire_87_43, c6288_wire_87_44, c6288_wire_87_45, c6288_wire_87_46});
fanout_n #(47, 0, 0) FANOUT_720 (c6288_wire_90, {c6288_wire_90_0, c6288_wire_90_1, c6288_wire_90_2, c6288_wire_90_3, c6288_wire_90_4, c6288_wire_90_5, c6288_wire_90_6, c6288_wire_90_7, c6288_wire_90_8, c6288_wire_90_9, c6288_wire_90_10, c6288_wire_90_11, c6288_wire_90_12, c6288_wire_90_13, c6288_wire_90_14, c6288_wire_90_15, c6288_wire_90_16, c6288_wire_90_17, c6288_wire_90_18, c6288_wire_90_19, c6288_wire_90_20, c6288_wire_90_21, c6288_wire_90_22, c6288_wire_90_23, c6288_wire_90_24, c6288_wire_90_25, c6288_wire_90_26, c6288_wire_90_27, c6288_wire_90_28, c6288_wire_90_29, c6288_wire_90_30, c6288_wire_90_31, c6288_wire_90_32, c6288_wire_90_33, c6288_wire_90_34, c6288_wire_90_35, c6288_wire_90_36, c6288_wire_90_37, c6288_wire_90_38, c6288_wire_90_39, c6288_wire_90_40, c6288_wire_90_41, c6288_wire_90_42, c6288_wire_90_43, c6288_wire_90_44, c6288_wire_90_45, c6288_wire_90_46});
fanout_n #(47, 0, 0) FANOUT_721 (c6288_wire_93, {c6288_wire_93_0, c6288_wire_93_1, c6288_wire_93_2, c6288_wire_93_3, c6288_wire_93_4, c6288_wire_93_5, c6288_wire_93_6, c6288_wire_93_7, c6288_wire_93_8, c6288_wire_93_9, c6288_wire_93_10, c6288_wire_93_11, c6288_wire_93_12, c6288_wire_93_13, c6288_wire_93_14, c6288_wire_93_15, c6288_wire_93_16, c6288_wire_93_17, c6288_wire_93_18, c6288_wire_93_19, c6288_wire_93_20, c6288_wire_93_21, c6288_wire_93_22, c6288_wire_93_23, c6288_wire_93_24, c6288_wire_93_25, c6288_wire_93_26, c6288_wire_93_27, c6288_wire_93_28, c6288_wire_93_29, c6288_wire_93_30, c6288_wire_93_31, c6288_wire_93_32, c6288_wire_93_33, c6288_wire_93_34, c6288_wire_93_35, c6288_wire_93_36, c6288_wire_93_37, c6288_wire_93_38, c6288_wire_93_39, c6288_wire_93_40, c6288_wire_93_41, c6288_wire_93_42, c6288_wire_93_43, c6288_wire_93_44, c6288_wire_93_45, c6288_wire_93_46});
fanout_n #(47, 0, 0) FANOUT_722 (c6288_wire_96, {c6288_wire_96_0, c6288_wire_96_1, c6288_wire_96_2, c6288_wire_96_3, c6288_wire_96_4, c6288_wire_96_5, c6288_wire_96_6, c6288_wire_96_7, c6288_wire_96_8, c6288_wire_96_9, c6288_wire_96_10, c6288_wire_96_11, c6288_wire_96_12, c6288_wire_96_13, c6288_wire_96_14, c6288_wire_96_15, c6288_wire_96_16, c6288_wire_96_17, c6288_wire_96_18, c6288_wire_96_19, c6288_wire_96_20, c6288_wire_96_21, c6288_wire_96_22, c6288_wire_96_23, c6288_wire_96_24, c6288_wire_96_25, c6288_wire_96_26, c6288_wire_96_27, c6288_wire_96_28, c6288_wire_96_29, c6288_wire_96_30, c6288_wire_96_31, c6288_wire_96_32, c6288_wire_96_33, c6288_wire_96_34, c6288_wire_96_35, c6288_wire_96_36, c6288_wire_96_37, c6288_wire_96_38, c6288_wire_96_39, c6288_wire_96_40, c6288_wire_96_41, c6288_wire_96_42, c6288_wire_96_43, c6288_wire_96_44, c6288_wire_96_45, c6288_wire_96_46});
fanout_n #(47, 0, 0) FANOUT_723 (c6288_wire_99, {c6288_wire_99_0, c6288_wire_99_1, c6288_wire_99_2, c6288_wire_99_3, c6288_wire_99_4, c6288_wire_99_5, c6288_wire_99_6, c6288_wire_99_7, c6288_wire_99_8, c6288_wire_99_9, c6288_wire_99_10, c6288_wire_99_11, c6288_wire_99_12, c6288_wire_99_13, c6288_wire_99_14, c6288_wire_99_15, c6288_wire_99_16, c6288_wire_99_17, c6288_wire_99_18, c6288_wire_99_19, c6288_wire_99_20, c6288_wire_99_21, c6288_wire_99_22, c6288_wire_99_23, c6288_wire_99_24, c6288_wire_99_25, c6288_wire_99_26, c6288_wire_99_27, c6288_wire_99_28, c6288_wire_99_29, c6288_wire_99_30, c6288_wire_99_31, c6288_wire_99_32, c6288_wire_99_33, c6288_wire_99_34, c6288_wire_99_35, c6288_wire_99_36, c6288_wire_99_37, c6288_wire_99_38, c6288_wire_99_39, c6288_wire_99_40, c6288_wire_99_41, c6288_wire_99_42, c6288_wire_99_43, c6288_wire_99_44, c6288_wire_99_45, c6288_wire_99_46});
fanout_n #(47, 0, 0) FANOUT_724 (c6288_wire_102, {c6288_wire_102_0, c6288_wire_102_1, c6288_wire_102_2, c6288_wire_102_3, c6288_wire_102_4, c6288_wire_102_5, c6288_wire_102_6, c6288_wire_102_7, c6288_wire_102_8, c6288_wire_102_9, c6288_wire_102_10, c6288_wire_102_11, c6288_wire_102_12, c6288_wire_102_13, c6288_wire_102_14, c6288_wire_102_15, c6288_wire_102_16, c6288_wire_102_17, c6288_wire_102_18, c6288_wire_102_19, c6288_wire_102_20, c6288_wire_102_21, c6288_wire_102_22, c6288_wire_102_23, c6288_wire_102_24, c6288_wire_102_25, c6288_wire_102_26, c6288_wire_102_27, c6288_wire_102_28, c6288_wire_102_29, c6288_wire_102_30, c6288_wire_102_31, c6288_wire_102_32, c6288_wire_102_33, c6288_wire_102_34, c6288_wire_102_35, c6288_wire_102_36, c6288_wire_102_37, c6288_wire_102_38, c6288_wire_102_39, c6288_wire_102_40, c6288_wire_102_41, c6288_wire_102_42, c6288_wire_102_43, c6288_wire_102_44, c6288_wire_102_45, c6288_wire_102_46});
fanout_n #(47, 0, 0) FANOUT_725 (c6288_wire_105, {c6288_wire_105_0, c6288_wire_105_1, c6288_wire_105_2, c6288_wire_105_3, c6288_wire_105_4, c6288_wire_105_5, c6288_wire_105_6, c6288_wire_105_7, c6288_wire_105_8, c6288_wire_105_9, c6288_wire_105_10, c6288_wire_105_11, c6288_wire_105_12, c6288_wire_105_13, c6288_wire_105_14, c6288_wire_105_15, c6288_wire_105_16, c6288_wire_105_17, c6288_wire_105_18, c6288_wire_105_19, c6288_wire_105_20, c6288_wire_105_21, c6288_wire_105_22, c6288_wire_105_23, c6288_wire_105_24, c6288_wire_105_25, c6288_wire_105_26, c6288_wire_105_27, c6288_wire_105_28, c6288_wire_105_29, c6288_wire_105_30, c6288_wire_105_31, c6288_wire_105_32, c6288_wire_105_33, c6288_wire_105_34, c6288_wire_105_35, c6288_wire_105_36, c6288_wire_105_37, c6288_wire_105_38, c6288_wire_105_39, c6288_wire_105_40, c6288_wire_105_41, c6288_wire_105_42, c6288_wire_105_43, c6288_wire_105_44, c6288_wire_105_45, c6288_wire_105_46});
fanout_n #(47, 0, 0) FANOUT_726 (c6288_wire_108, {c6288_wire_108_0, c6288_wire_108_1, c6288_wire_108_2, c6288_wire_108_3, c6288_wire_108_4, c6288_wire_108_5, c6288_wire_108_6, c6288_wire_108_7, c6288_wire_108_8, c6288_wire_108_9, c6288_wire_108_10, c6288_wire_108_11, c6288_wire_108_12, c6288_wire_108_13, c6288_wire_108_14, c6288_wire_108_15, c6288_wire_108_16, c6288_wire_108_17, c6288_wire_108_18, c6288_wire_108_19, c6288_wire_108_20, c6288_wire_108_21, c6288_wire_108_22, c6288_wire_108_23, c6288_wire_108_24, c6288_wire_108_25, c6288_wire_108_26, c6288_wire_108_27, c6288_wire_108_28, c6288_wire_108_29, c6288_wire_108_30, c6288_wire_108_31, c6288_wire_108_32, c6288_wire_108_33, c6288_wire_108_34, c6288_wire_108_35, c6288_wire_108_36, c6288_wire_108_37, c6288_wire_108_38, c6288_wire_108_39, c6288_wire_108_40, c6288_wire_108_41, c6288_wire_108_42, c6288_wire_108_43, c6288_wire_108_44, c6288_wire_108_45, c6288_wire_108_46});
fanout_n #(47, 0, 0) FANOUT_727 (c6288_wire_111, {c6288_wire_111_0, c6288_wire_111_1, c6288_wire_111_2, c6288_wire_111_3, c6288_wire_111_4, c6288_wire_111_5, c6288_wire_111_6, c6288_wire_111_7, c6288_wire_111_8, c6288_wire_111_9, c6288_wire_111_10, c6288_wire_111_11, c6288_wire_111_12, c6288_wire_111_13, c6288_wire_111_14, c6288_wire_111_15, c6288_wire_111_16, c6288_wire_111_17, c6288_wire_111_18, c6288_wire_111_19, c6288_wire_111_20, c6288_wire_111_21, c6288_wire_111_22, c6288_wire_111_23, c6288_wire_111_24, c6288_wire_111_25, c6288_wire_111_26, c6288_wire_111_27, c6288_wire_111_28, c6288_wire_111_29, c6288_wire_111_30, c6288_wire_111_31, c6288_wire_111_32, c6288_wire_111_33, c6288_wire_111_34, c6288_wire_111_35, c6288_wire_111_36, c6288_wire_111_37, c6288_wire_111_38, c6288_wire_111_39, c6288_wire_111_40, c6288_wire_111_41, c6288_wire_111_42, c6288_wire_111_43, c6288_wire_111_44, c6288_wire_111_45, c6288_wire_111_46});
fanout_n #(47, 0, 0) FANOUT_728 (c6288_wire_114, {c6288_wire_114_0, c6288_wire_114_1, c6288_wire_114_2, c6288_wire_114_3, c6288_wire_114_4, c6288_wire_114_5, c6288_wire_114_6, c6288_wire_114_7, c6288_wire_114_8, c6288_wire_114_9, c6288_wire_114_10, c6288_wire_114_11, c6288_wire_114_12, c6288_wire_114_13, c6288_wire_114_14, c6288_wire_114_15, c6288_wire_114_16, c6288_wire_114_17, c6288_wire_114_18, c6288_wire_114_19, c6288_wire_114_20, c6288_wire_114_21, c6288_wire_114_22, c6288_wire_114_23, c6288_wire_114_24, c6288_wire_114_25, c6288_wire_114_26, c6288_wire_114_27, c6288_wire_114_28, c6288_wire_114_29, c6288_wire_114_30, c6288_wire_114_31, c6288_wire_114_32, c6288_wire_114_33, c6288_wire_114_34, c6288_wire_114_35, c6288_wire_114_36, c6288_wire_114_37, c6288_wire_114_38, c6288_wire_114_39, c6288_wire_114_40, c6288_wire_114_41, c6288_wire_114_42, c6288_wire_114_43, c6288_wire_114_44, c6288_wire_114_45, c6288_wire_114_46});
fanout_n #(46, 0, 0) FANOUT_729 (c6288_wire_42, {c6288_wire_42_0, c6288_wire_42_1, c6288_wire_42_2, c6288_wire_42_3, c6288_wire_42_4, c6288_wire_42_5, c6288_wire_42_6, c6288_wire_42_7, c6288_wire_42_8, c6288_wire_42_9, c6288_wire_42_10, c6288_wire_42_11, c6288_wire_42_12, c6288_wire_42_13, c6288_wire_42_14, c6288_wire_42_15, c6288_wire_42_16, c6288_wire_42_17, c6288_wire_42_18, c6288_wire_42_19, c6288_wire_42_20, c6288_wire_42_21, c6288_wire_42_22, c6288_wire_42_23, c6288_wire_42_24, c6288_wire_42_25, c6288_wire_42_26, c6288_wire_42_27, c6288_wire_42_28, c6288_wire_42_29, c6288_wire_42_30, c6288_wire_42_31, c6288_wire_42_32, c6288_wire_42_33, c6288_wire_42_34, c6288_wire_42_35, c6288_wire_42_36, c6288_wire_42_37, c6288_wire_42_38, c6288_wire_42_39, c6288_wire_42_40, c6288_wire_42_41, c6288_wire_42_42, c6288_wire_42_43, c6288_wire_42_44, c6288_wire_42_45});
fanout_n #(47, 0, 0) FANOUT_730 (c6288_wire_117, {c6288_wire_117_0, c6288_wire_117_1, c6288_wire_117_2, c6288_wire_117_3, c6288_wire_117_4, c6288_wire_117_5, c6288_wire_117_6, c6288_wire_117_7, c6288_wire_117_8, c6288_wire_117_9, c6288_wire_117_10, c6288_wire_117_11, c6288_wire_117_12, c6288_wire_117_13, c6288_wire_117_14, c6288_wire_117_15, c6288_wire_117_16, c6288_wire_117_17, c6288_wire_117_18, c6288_wire_117_19, c6288_wire_117_20, c6288_wire_117_21, c6288_wire_117_22, c6288_wire_117_23, c6288_wire_117_24, c6288_wire_117_25, c6288_wire_117_26, c6288_wire_117_27, c6288_wire_117_28, c6288_wire_117_29, c6288_wire_117_30, c6288_wire_117_31, c6288_wire_117_32, c6288_wire_117_33, c6288_wire_117_34, c6288_wire_117_35, c6288_wire_117_36, c6288_wire_117_37, c6288_wire_117_38, c6288_wire_117_39, c6288_wire_117_40, c6288_wire_117_41, c6288_wire_117_42, c6288_wire_117_43, c6288_wire_117_44, c6288_wire_117_45, c6288_wire_117_46});
fanout_n #(46, 0, 0) FANOUT_731 (c6288_wire_47, {c6288_wire_47_0, c6288_wire_47_1, c6288_wire_47_2, c6288_wire_47_3, c6288_wire_47_4, c6288_wire_47_5, c6288_wire_47_6, c6288_wire_47_7, c6288_wire_47_8, c6288_wire_47_9, c6288_wire_47_10, c6288_wire_47_11, c6288_wire_47_12, c6288_wire_47_13, c6288_wire_47_14, c6288_wire_47_15, c6288_wire_47_16, c6288_wire_47_17, c6288_wire_47_18, c6288_wire_47_19, c6288_wire_47_20, c6288_wire_47_21, c6288_wire_47_22, c6288_wire_47_23, c6288_wire_47_24, c6288_wire_47_25, c6288_wire_47_26, c6288_wire_47_27, c6288_wire_47_28, c6288_wire_47_29, c6288_wire_47_30, c6288_wire_47_31, c6288_wire_47_32, c6288_wire_47_33, c6288_wire_47_34, c6288_wire_47_35, c6288_wire_47_36, c6288_wire_47_37, c6288_wire_47_38, c6288_wire_47_39, c6288_wire_47_40, c6288_wire_47_41, c6288_wire_47_42, c6288_wire_47_43, c6288_wire_47_44, c6288_wire_47_45});
fanout_n #(46, 0, 0) FANOUT_732 (c6288_wire_52, {c6288_wire_52_0, c6288_wire_52_1, c6288_wire_52_2, c6288_wire_52_3, c6288_wire_52_4, c6288_wire_52_5, c6288_wire_52_6, c6288_wire_52_7, c6288_wire_52_8, c6288_wire_52_9, c6288_wire_52_10, c6288_wire_52_11, c6288_wire_52_12, c6288_wire_52_13, c6288_wire_52_14, c6288_wire_52_15, c6288_wire_52_16, c6288_wire_52_17, c6288_wire_52_18, c6288_wire_52_19, c6288_wire_52_20, c6288_wire_52_21, c6288_wire_52_22, c6288_wire_52_23, c6288_wire_52_24, c6288_wire_52_25, c6288_wire_52_26, c6288_wire_52_27, c6288_wire_52_28, c6288_wire_52_29, c6288_wire_52_30, c6288_wire_52_31, c6288_wire_52_32, c6288_wire_52_33, c6288_wire_52_34, c6288_wire_52_35, c6288_wire_52_36, c6288_wire_52_37, c6288_wire_52_38, c6288_wire_52_39, c6288_wire_52_40, c6288_wire_52_41, c6288_wire_52_42, c6288_wire_52_43, c6288_wire_52_44, c6288_wire_52_45});


and_n #(2, 0, 0) AND_1 (c6288_wire_1, {c6288_wire_2_0, c6288_wire_3_0});
and_n #(3, 0, 0) AND_2 (c6288_wire_4, {c6288_wire_1_0, c6288_wire_5_0, c6288_wire_6_0});
notg #(0, 0) NOT_1 (c6288_wire_7, c6288_wire_1_1);
and_n #(3, 0, 0) AND_3 (c6288_wire_8, {c6288_wire_1_2, c6288_wire_5_1, c6288_wire_6_1});
and_n #(2, 0, 0) AND_4 (c6288_wire_9, {c6288_wire_10_0, c6288_wire_3_1});
and_n #(3, 0, 0) AND_5 (c6288_wire_11, {c6288_wire_9_0, c6288_wire_2_1, c6288_wire_6_2});
notg #(0, 0) NOT_2 (c6288_wire_12, c6288_wire_9_1);
and_n #(3, 0, 0) AND_6 (c6288_wire_13, {c6288_wire_9_2, c6288_wire_2_2, c6288_wire_6_3});
and_n #(2, 0, 0) AND_7 (c6288_wire_14, {c6288_wire_15_0, c6288_wire_3_2});
and_n #(3, 0, 0) AND_8 (c6288_wire_16, {c6288_wire_14_0, c6288_wire_10_1, c6288_wire_6_4});
notg #(0, 0) NOT_3 (c6288_wire_17, c6288_wire_14_1);
and_n #(3, 0, 0) AND_9 (c6288_wire_18, {c6288_wire_14_2, c6288_wire_10_2, c6288_wire_6_5});
and_n #(2, 0, 0) AND_10 (c6288_wire_19, {c6288_wire_20_0, c6288_wire_3_3});
and_n #(3, 0, 0) AND_11 (c6288_wire_21, {c6288_wire_19_0, c6288_wire_15_1, c6288_wire_6_6});
notg #(0, 0) NOT_4 (c6288_wire_22, c6288_wire_19_1);
and_n #(3, 0, 0) AND_12 (c6288_wire_23, {c6288_wire_19_2, c6288_wire_15_2, c6288_wire_6_7});
and_n #(2, 0, 0) AND_13 (c6288_wire_24, {c6288_wire_25_0, c6288_wire_3_4});
and_n #(3, 0, 0) AND_14 (c6288_wire_26, {c6288_wire_24_0, c6288_wire_20_1, c6288_wire_6_8});
notg #(0, 0) NOT_5 (c6288_wire_27, c6288_wire_24_1);
and_n #(3, 0, 0) AND_15 (c6288_wire_28, {c6288_wire_24_2, c6288_wire_20_2, c6288_wire_6_9});
and_n #(2, 0, 0) AND_16 (c6288_wire_29, {c6288_wire_30_0, c6288_wire_3_5});
and_n #(3, 0, 0) AND_17 (c6288_wire_31, {c6288_wire_29_0, c6288_wire_32_0, c6288_wire_6_10});
notg #(0, 0) NOT_6 (c6288_wire_33, c6288_wire_29_1);
and_n #(2, 0, 0) AND_18 (c6288_wire_34, {c6288_wire_29_2, c6288_wire_35});
and_n #(2, 0, 0) AND_19 (c6288_wire_36, {c6288_wire_37_0, c6288_wire_3_6});
and_n #(3, 0, 0) AND_20 (c6288_wire_38, {c6288_wire_36_0, c6288_wire_30_1, c6288_wire_6_11});
notg #(0, 0) NOT_7 (c6288_wire_39, c6288_wire_36_1);
and_n #(3, 0, 0) AND_21 (c6288_wire_40, {c6288_wire_36_2, c6288_wire_30_2, c6288_wire_6_12});
and_n #(2, 0, 0) AND_22 (c6288_wire_41, {c6288_wire_42_0, c6288_wire_3_7});
and_n #(3, 0, 0) AND_23 (c6288_wire_43, {c6288_wire_41_0, c6288_wire_37_1, c6288_wire_6_13});
notg #(0, 0) NOT_8 (c6288_wire_44, c6288_wire_41_1);
and_n #(3, 0, 0) AND_24 (c6288_wire_45, {c6288_wire_41_2, c6288_wire_37_2, c6288_wire_6_14});
and_n #(2, 0, 0) AND_25 (c6288_wire_46, {c6288_wire_47_0, c6288_wire_3_8});
and_n #(3, 0, 0) AND_26 (c6288_wire_48, {c6288_wire_46_0, c6288_wire_42_1, c6288_wire_6_15});
notg #(0, 0) NOT_9 (c6288_wire_49, c6288_wire_46_1);
and_n #(3, 0, 0) AND_27 (c6288_wire_50, {c6288_wire_46_2, c6288_wire_42_2, c6288_wire_6_16});
and_n #(2, 0, 0) AND_28 (c6288_wire_51, {c6288_wire_52_0, c6288_wire_3_9});
and_n #(3, 0, 0) AND_29 (c6288_wire_53, {c6288_wire_51_0, c6288_wire_47_1, c6288_wire_6_17});
notg #(0, 0) NOT_10 (c6288_wire_54, c6288_wire_51_1);
and_n #(3, 0, 0) AND_30 (c6288_wire_55, {c6288_wire_51_2, c6288_wire_47_2, c6288_wire_6_18});
and_n #(2, 0, 0) AND_31 (c6288_wire_56, {c6288_wire_57_0, c6288_wire_3_10});
and_n #(3, 0, 0) AND_32 (c6288_wire_58, {c6288_wire_56_0, c6288_wire_52_1, c6288_wire_6_19});
notg #(0, 0) NOT_11 (c6288_wire_59, c6288_wire_56_1);
and_n #(3, 0, 0) AND_33 (c6288_wire_60, {c6288_wire_56_2, c6288_wire_52_2, c6288_wire_6_20});
and_n #(2, 0, 0) AND_34 (c6288_wire_61, {c6288_wire_62_0, c6288_wire_3_11});
and_n #(3, 0, 0) AND_35 (c6288_wire_63, {c6288_wire_61_0, c6288_wire_57_1, c6288_wire_6_21});
notg #(0, 0) NOT_12 (c6288_wire_64, c6288_wire_61_1);
and_n #(3, 0, 0) AND_36 (c6288_wire_65, {c6288_wire_61_2, c6288_wire_57_2, c6288_wire_6_22});
and_n #(2, 0, 0) AND_37 (c6288_wire_66, {c6288_wire_67_0, c6288_wire_3_12});
and_n #(3, 0, 0) AND_38 (c6288_wire_68, {c6288_wire_66_0, c6288_wire_62_1, c6288_wire_6_23});
notg #(0, 0) NOT_13 (c6288_wire_69, c6288_wire_66_1);
and_n #(3, 0, 0) AND_39 (c6288_wire_70, {c6288_wire_66_2, c6288_wire_62_2, c6288_wire_6_24});
and_n #(2, 0, 0) AND_40 (c6288_wire_71, {c6288_wire_5_2, c6288_wire_3_13});
and_n #(3, 0, 0) AND_41 (c6288_wire_72, {c6288_wire_71_0, c6288_wire_67_1, c6288_wire_6_25});
notg #(0, 0) NOT_14 (c6288_wire_73, c6288_wire_71_1);
and_n #(3, 0, 0) AND_42 (c6288_wire_74, {c6288_wire_71_2, c6288_wire_67_2, c6288_wire_6_26});
and_n #(2, 0, 0) AND_43 (c6288_wire_75, {c6288_wire_32_1, c6288_wire_3_14});
and_n #(2, 0, 0) AND_44 (c6288_wire_76, {c6288_wire_32_2, c6288_wire_6_27});
and_n #(2, 0, 0) AND_45 (c6288_wire_77, {c6288_wire_32_3, c6288_wire_78_0});
and_n #(2, 0, 0) AND_46 (c6288_wire_79, {c6288_wire_32_4, c6288_wire_78_1});
and_n #(2, 0, 0) AND_47 (c6288_wire_80, {c6288_wire_32_5, c6288_wire_81_0});
and_n #(2, 0, 0) AND_48 (c6288_wire_82, {c6288_wire_32_6, c6288_wire_81_1});
and_n #(2, 0, 0) AND_49 (c6288_wire_83, {c6288_wire_32_7, c6288_wire_84_0});
and_n #(2, 0, 0) AND_50 (c6288_wire_85, {c6288_wire_32_8, c6288_wire_84_1});
and_n #(2, 0, 0) AND_51 (c6288_wire_86, {c6288_wire_32_9, c6288_wire_87_0});
and_n #(2, 0, 0) AND_52 (c6288_wire_88, {c6288_wire_32_10, c6288_wire_87_1});
and_n #(2, 0, 0) AND_53 (c6288_wire_89, {c6288_wire_32_11, c6288_wire_90_0});
and_n #(2, 0, 0) AND_54 (c6288_wire_91, {c6288_wire_32_12, c6288_wire_90_1});
and_n #(2, 0, 0) AND_55 (c6288_wire_92, {c6288_wire_32_13, c6288_wire_93_0});
and_n #(2, 0, 0) AND_56 (c6288_wire_94, {c6288_wire_32_14, c6288_wire_93_1});
and_n #(2, 0, 0) AND_57 (c6288_wire_95, {c6288_wire_32_15, c6288_wire_96_0});
and_n #(2, 0, 0) AND_58 (c6288_wire_97, {c6288_wire_32_16, c6288_wire_96_1});
and_n #(2, 0, 0) AND_59 (c6288_wire_98, {c6288_wire_32_17, c6288_wire_99_0});
and_n #(2, 0, 0) AND_60 (c6288_wire_100, {c6288_wire_32_18, c6288_wire_99_1});
and_n #(2, 0, 0) AND_61 (c6288_wire_101, {c6288_wire_32_19, c6288_wire_102_0});
and_n #(2, 0, 0) AND_62 (c6288_wire_103, {c6288_wire_32_20, c6288_wire_102_1});
and_n #(2, 0, 0) AND_63 (c6288_wire_104, {c6288_wire_32_21, c6288_wire_105_0});
and_n #(2, 0, 0) AND_64 (c6288_wire_106, {c6288_wire_32_22, c6288_wire_105_1});
and_n #(2, 0, 0) AND_65 (c6288_wire_107, {c6288_wire_32_23, c6288_wire_108_0});
and_n #(2, 0, 0) AND_66 (c6288_wire_109, {c6288_wire_32_24, c6288_wire_108_1});
and_n #(2, 0, 0) AND_67 (c6288_wire_110, {c6288_wire_32_25, c6288_wire_111_0});
and_n #(2, 0, 0) AND_68 (c6288_wire_112, {c6288_wire_32_26, c6288_wire_111_1});
and_n #(2, 0, 0) AND_69 (c6288_wire_113, {c6288_wire_32_27, c6288_wire_114_0});
and_n #(2, 0, 0) AND_70 (c6288_wire_115, {c6288_wire_32_28, c6288_wire_114_1});
and_n #(2, 0, 0) AND_71 (c6288_wire_116, {c6288_wire_32_29, c6288_wire_117_0});
and_n #(2, 0, 0) AND_72 (c6288_wire_118, {c6288_wire_32_30, c6288_wire_117_1});
and_n #(2, 0, 0) AND_73 (c6288_wire_119, {c6288_wire_2_3, c6288_wire_78_2});
and_n #(2, 0, 0) AND_74 (c6288_wire_120, {c6288_wire_2_4, c6288_wire_81_2});
and_n #(2, 0, 0) AND_75 (c6288_wire_121, {c6288_wire_2_5, c6288_wire_84_2});
and_n #(2, 0, 0) AND_76 (c6288_wire_122, {c6288_wire_2_6, c6288_wire_87_2});
and_n #(2, 0, 0) AND_77 (c6288_wire_123, {c6288_wire_2_7, c6288_wire_90_2});
and_n #(2, 0, 0) AND_78 (c6288_wire_124, {c6288_wire_2_8, c6288_wire_93_2});
and_n #(2, 0, 0) AND_79 (c6288_wire_125, {c6288_wire_2_9, c6288_wire_96_2});
and_n #(2, 0, 0) AND_80 (c6288_wire_126, {c6288_wire_2_10, c6288_wire_99_2});
and_n #(2, 0, 0) AND_81 (c6288_wire_127, {c6288_wire_2_11, c6288_wire_102_2});
and_n #(2, 0, 0) AND_82 (c6288_wire_128, {c6288_wire_2_12, c6288_wire_105_2});
and_n #(2, 0, 0) AND_83 (c6288_wire_129, {c6288_wire_2_13, c6288_wire_108_2});
and_n #(2, 0, 0) AND_84 (c6288_wire_130, {c6288_wire_2_14, c6288_wire_111_2});
and_n #(2, 0, 0) AND_85 (c6288_wire_131, {c6288_wire_2_15, c6288_wire_114_2});
and_n #(2, 0, 0) AND_86 (c6288_wire_132, {c6288_wire_2_16, c6288_wire_117_2});
and_n #(3, 0, 0) AND_87 (c6288_wire_133, {c6288_wire_2_17, c6288_wire_117_3, c6288_wire_134_0});
and_n #(3, 0, 0) AND_88 (c6288_wire_135, {c6288_wire_2_18, c6288_wire_114_3, c6288_wire_136_0});
and_n #(3, 0, 0) AND_89 (c6288_wire_137, {c6288_wire_2_19, c6288_wire_111_3, c6288_wire_138_0});
and_n #(3, 0, 0) AND_90 (c6288_wire_139, {c6288_wire_2_20, c6288_wire_108_3, c6288_wire_140_0});
and_n #(3, 0, 0) AND_91 (c6288_wire_141, {c6288_wire_2_21, c6288_wire_105_3, c6288_wire_142_0});
and_n #(3, 0, 0) AND_92 (c6288_wire_143, {c6288_wire_2_22, c6288_wire_102_3, c6288_wire_144_0});
and_n #(3, 0, 0) AND_93 (c6288_wire_145, {c6288_wire_2_23, c6288_wire_99_3, c6288_wire_146_0});
and_n #(3, 0, 0) AND_94 (c6288_wire_147, {c6288_wire_2_24, c6288_wire_96_3, c6288_wire_148_0});
and_n #(3, 0, 0) AND_95 (c6288_wire_149, {c6288_wire_2_25, c6288_wire_93_3, c6288_wire_150_0});
and_n #(3, 0, 0) AND_96 (c6288_wire_151, {c6288_wire_2_26, c6288_wire_90_3, c6288_wire_152_0});
and_n #(3, 0, 0) AND_97 (c6288_wire_153, {c6288_wire_2_27, c6288_wire_87_3, c6288_wire_154_0});
and_n #(3, 0, 0) AND_98 (c6288_wire_155, {c6288_wire_2_28, c6288_wire_84_3, c6288_wire_156_0});
and_n #(3, 0, 0) AND_99 (c6288_wire_157, {c6288_wire_2_29, c6288_wire_81_3, c6288_wire_158_0});
and_n #(3, 0, 0) AND_100 (c6288_wire_159, {c6288_wire_2_30, c6288_wire_78_3, c6288_wire_160_0});
and_n #(2, 0, 0) AND_101 (c6288_wire_161, {c6288_wire_10_3, c6288_wire_78_4});
and_n #(2, 0, 0) AND_102 (c6288_wire_162, {c6288_wire_10_4, c6288_wire_81_4});
and_n #(2, 0, 0) AND_103 (c6288_wire_163, {c6288_wire_10_5, c6288_wire_84_4});
and_n #(2, 0, 0) AND_104 (c6288_wire_164, {c6288_wire_10_6, c6288_wire_87_4});
and_n #(2, 0, 0) AND_105 (c6288_wire_165, {c6288_wire_10_7, c6288_wire_90_4});
and_n #(2, 0, 0) AND_106 (c6288_wire_166, {c6288_wire_10_8, c6288_wire_93_4});
and_n #(2, 0, 0) AND_107 (c6288_wire_167, {c6288_wire_10_9, c6288_wire_96_4});
and_n #(2, 0, 0) AND_108 (c6288_wire_168, {c6288_wire_10_10, c6288_wire_99_4});
and_n #(2, 0, 0) AND_109 (c6288_wire_169, {c6288_wire_10_11, c6288_wire_102_4});
and_n #(2, 0, 0) AND_110 (c6288_wire_170, {c6288_wire_10_12, c6288_wire_105_4});
and_n #(2, 0, 0) AND_111 (c6288_wire_171, {c6288_wire_10_13, c6288_wire_108_4});
and_n #(2, 0, 0) AND_112 (c6288_wire_172, {c6288_wire_10_14, c6288_wire_111_4});
and_n #(2, 0, 0) AND_113 (c6288_wire_173, {c6288_wire_10_15, c6288_wire_114_4});
and_n #(2, 0, 0) AND_114 (c6288_wire_174, {c6288_wire_10_16, c6288_wire_117_4});
and_n #(3, 0, 0) AND_115 (c6288_wire_175, {c6288_wire_10_17, c6288_wire_117_5, c6288_wire_176_0});
and_n #(3, 0, 0) AND_116 (c6288_wire_177, {c6288_wire_10_18, c6288_wire_114_5, c6288_wire_178_0});
and_n #(3, 0, 0) AND_117 (c6288_wire_179, {c6288_wire_10_19, c6288_wire_111_5, c6288_wire_180_0});
and_n #(3, 0, 0) AND_118 (c6288_wire_181, {c6288_wire_10_20, c6288_wire_108_5, c6288_wire_182_0});
and_n #(3, 0, 0) AND_119 (c6288_wire_183, {c6288_wire_10_21, c6288_wire_105_5, c6288_wire_184_0});
and_n #(3, 0, 0) AND_120 (c6288_wire_185, {c6288_wire_10_22, c6288_wire_102_5, c6288_wire_186_0});
and_n #(3, 0, 0) AND_121 (c6288_wire_187, {c6288_wire_10_23, c6288_wire_99_5, c6288_wire_188_0});
and_n #(3, 0, 0) AND_122 (c6288_wire_189, {c6288_wire_10_24, c6288_wire_96_5, c6288_wire_190_0});
and_n #(3, 0, 0) AND_123 (c6288_wire_191, {c6288_wire_10_25, c6288_wire_93_5, c6288_wire_192_0});
and_n #(3, 0, 0) AND_124 (c6288_wire_193, {c6288_wire_10_26, c6288_wire_90_5, c6288_wire_194_0});
and_n #(3, 0, 0) AND_125 (c6288_wire_195, {c6288_wire_10_27, c6288_wire_87_5, c6288_wire_196_0});
and_n #(3, 0, 0) AND_126 (c6288_wire_197, {c6288_wire_10_28, c6288_wire_84_5, c6288_wire_198_0});
and_n #(3, 0, 0) AND_127 (c6288_wire_199, {c6288_wire_10_29, c6288_wire_81_5, c6288_wire_200_0});
and_n #(3, 0, 0) AND_128 (c6288_wire_201, {c6288_wire_10_30, c6288_wire_78_5, c6288_wire_202_0});
and_n #(2, 0, 0) AND_129 (c6288_wire_203, {c6288_wire_15_3, c6288_wire_78_6});
and_n #(2, 0, 0) AND_130 (c6288_wire_204, {c6288_wire_15_4, c6288_wire_81_6});
and_n #(2, 0, 0) AND_131 (c6288_wire_205, {c6288_wire_15_5, c6288_wire_84_6});
and_n #(2, 0, 0) AND_132 (c6288_wire_206, {c6288_wire_15_6, c6288_wire_87_6});
and_n #(2, 0, 0) AND_133 (c6288_wire_207, {c6288_wire_15_7, c6288_wire_90_6});
and_n #(2, 0, 0) AND_134 (c6288_wire_208, {c6288_wire_15_8, c6288_wire_93_6});
and_n #(2, 0, 0) AND_135 (c6288_wire_209, {c6288_wire_15_9, c6288_wire_96_6});
and_n #(2, 0, 0) AND_136 (c6288_wire_210, {c6288_wire_15_10, c6288_wire_99_6});
and_n #(2, 0, 0) AND_137 (c6288_wire_211, {c6288_wire_15_11, c6288_wire_102_6});
and_n #(2, 0, 0) AND_138 (c6288_wire_212, {c6288_wire_15_12, c6288_wire_105_6});
and_n #(2, 0, 0) AND_139 (c6288_wire_213, {c6288_wire_15_13, c6288_wire_108_6});
and_n #(2, 0, 0) AND_140 (c6288_wire_214, {c6288_wire_15_14, c6288_wire_111_6});
and_n #(2, 0, 0) AND_141 (c6288_wire_215, {c6288_wire_15_15, c6288_wire_114_6});
and_n #(2, 0, 0) AND_142 (c6288_wire_216, {c6288_wire_15_16, c6288_wire_117_6});
and_n #(3, 0, 0) AND_143 (c6288_wire_217, {c6288_wire_15_17, c6288_wire_117_7, c6288_wire_218_0});
and_n #(3, 0, 0) AND_144 (c6288_wire_219, {c6288_wire_15_18, c6288_wire_114_7, c6288_wire_220_0});
and_n #(3, 0, 0) AND_145 (c6288_wire_221, {c6288_wire_15_19, c6288_wire_111_7, c6288_wire_222_0});
and_n #(3, 0, 0) AND_146 (c6288_wire_223, {c6288_wire_15_20, c6288_wire_108_7, c6288_wire_224_0});
and_n #(3, 0, 0) AND_147 (c6288_wire_225, {c6288_wire_15_21, c6288_wire_105_7, c6288_wire_226_0});
and_n #(3, 0, 0) AND_148 (c6288_wire_227, {c6288_wire_15_22, c6288_wire_102_7, c6288_wire_228_0});
and_n #(3, 0, 0) AND_149 (c6288_wire_229, {c6288_wire_15_23, c6288_wire_99_7, c6288_wire_230_0});
and_n #(3, 0, 0) AND_150 (c6288_wire_231, {c6288_wire_15_24, c6288_wire_96_7, c6288_wire_232_0});
and_n #(3, 0, 0) AND_151 (c6288_wire_233, {c6288_wire_15_25, c6288_wire_93_7, c6288_wire_234_0});
and_n #(3, 0, 0) AND_152 (c6288_wire_235, {c6288_wire_15_26, c6288_wire_90_7, c6288_wire_236_0});
and_n #(3, 0, 0) AND_153 (c6288_wire_237, {c6288_wire_15_27, c6288_wire_87_7, c6288_wire_238_0});
and_n #(3, 0, 0) AND_154 (c6288_wire_239, {c6288_wire_15_28, c6288_wire_84_7, c6288_wire_240_0});
and_n #(3, 0, 0) AND_155 (c6288_wire_241, {c6288_wire_15_29, c6288_wire_81_7, c6288_wire_242_0});
and_n #(3, 0, 0) AND_156 (c6288_wire_243, {c6288_wire_15_30, c6288_wire_78_7, c6288_wire_244_0});
and_n #(2, 0, 0) AND_157 (c6288_wire_245, {c6288_wire_20_3, c6288_wire_78_8});
and_n #(2, 0, 0) AND_158 (c6288_wire_246, {c6288_wire_20_4, c6288_wire_81_8});
and_n #(2, 0, 0) AND_159 (c6288_wire_247, {c6288_wire_20_5, c6288_wire_84_8});
and_n #(2, 0, 0) AND_160 (c6288_wire_248, {c6288_wire_20_6, c6288_wire_87_8});
and_n #(2, 0, 0) AND_161 (c6288_wire_249, {c6288_wire_20_7, c6288_wire_90_8});
and_n #(2, 0, 0) AND_162 (c6288_wire_250, {c6288_wire_20_8, c6288_wire_93_8});
and_n #(2, 0, 0) AND_163 (c6288_wire_251, {c6288_wire_20_9, c6288_wire_96_8});
and_n #(2, 0, 0) AND_164 (c6288_wire_252, {c6288_wire_20_10, c6288_wire_99_8});
and_n #(2, 0, 0) AND_165 (c6288_wire_253, {c6288_wire_20_11, c6288_wire_102_8});
and_n #(2, 0, 0) AND_166 (c6288_wire_254, {c6288_wire_20_12, c6288_wire_105_8});
and_n #(2, 0, 0) AND_167 (c6288_wire_255, {c6288_wire_20_13, c6288_wire_108_8});
and_n #(2, 0, 0) AND_168 (c6288_wire_256, {c6288_wire_20_14, c6288_wire_111_8});
and_n #(2, 0, 0) AND_169 (c6288_wire_257, {c6288_wire_20_15, c6288_wire_114_8});
and_n #(2, 0, 0) AND_170 (c6288_wire_258, {c6288_wire_20_16, c6288_wire_117_8});
and_n #(3, 0, 0) AND_171 (c6288_wire_259, {c6288_wire_20_17, c6288_wire_117_9, c6288_wire_260_0});
and_n #(3, 0, 0) AND_172 (c6288_wire_261, {c6288_wire_20_18, c6288_wire_114_9, c6288_wire_262_0});
and_n #(3, 0, 0) AND_173 (c6288_wire_263, {c6288_wire_20_19, c6288_wire_111_9, c6288_wire_264_0});
and_n #(3, 0, 0) AND_174 (c6288_wire_265, {c6288_wire_20_20, c6288_wire_108_9, c6288_wire_266_0});
and_n #(3, 0, 0) AND_175 (c6288_wire_267, {c6288_wire_20_21, c6288_wire_105_9, c6288_wire_268_0});
and_n #(3, 0, 0) AND_176 (c6288_wire_269, {c6288_wire_20_22, c6288_wire_102_9, c6288_wire_270_0});
and_n #(3, 0, 0) AND_177 (c6288_wire_271, {c6288_wire_20_23, c6288_wire_99_9, c6288_wire_272_0});
and_n #(3, 0, 0) AND_178 (c6288_wire_273, {c6288_wire_20_24, c6288_wire_96_9, c6288_wire_274_0});
and_n #(3, 0, 0) AND_179 (c6288_wire_275, {c6288_wire_20_25, c6288_wire_93_9, c6288_wire_276_0});
and_n #(3, 0, 0) AND_180 (c6288_wire_277, {c6288_wire_20_26, c6288_wire_90_9, c6288_wire_278_0});
and_n #(3, 0, 0) AND_181 (c6288_wire_279, {c6288_wire_20_27, c6288_wire_87_9, c6288_wire_280_0});
and_n #(3, 0, 0) AND_182 (c6288_wire_281, {c6288_wire_20_28, c6288_wire_84_9, c6288_wire_282_0});
and_n #(3, 0, 0) AND_183 (c6288_wire_283, {c6288_wire_20_29, c6288_wire_81_9, c6288_wire_284_0});
and_n #(3, 0, 0) AND_184 (c6288_wire_285, {c6288_wire_20_30, c6288_wire_78_9, c6288_wire_286_0});
and_n #(2, 0, 0) AND_185 (c6288_wire_287, {c6288_wire_25_1, c6288_wire_78_10});
and_n #(2, 0, 0) AND_186 (c6288_wire_288, {c6288_wire_25_2, c6288_wire_78_11});
and_n #(2, 0, 0) AND_187 (c6288_wire_289, {c6288_wire_25_3, c6288_wire_81_10});
and_n #(2, 0, 0) AND_188 (c6288_wire_290, {c6288_wire_25_4, c6288_wire_84_10});
and_n #(2, 0, 0) AND_189 (c6288_wire_291, {c6288_wire_25_5, c6288_wire_87_10});
and_n #(2, 0, 0) AND_190 (c6288_wire_292, {c6288_wire_25_6, c6288_wire_90_10});
and_n #(2, 0, 0) AND_191 (c6288_wire_293, {c6288_wire_25_7, c6288_wire_93_10});
and_n #(2, 0, 0) AND_192 (c6288_wire_294, {c6288_wire_25_8, c6288_wire_96_10});
and_n #(2, 0, 0) AND_193 (c6288_wire_295, {c6288_wire_25_9, c6288_wire_99_10});
and_n #(2, 0, 0) AND_194 (c6288_wire_296, {c6288_wire_25_10, c6288_wire_102_10});
and_n #(2, 0, 0) AND_195 (c6288_wire_297, {c6288_wire_25_11, c6288_wire_105_10});
and_n #(2, 0, 0) AND_196 (c6288_wire_298, {c6288_wire_25_12, c6288_wire_108_10});
and_n #(2, 0, 0) AND_197 (c6288_wire_299, {c6288_wire_25_13, c6288_wire_111_10});
and_n #(2, 0, 0) AND_198 (c6288_wire_300, {c6288_wire_25_14, c6288_wire_114_10});
and_n #(2, 0, 0) AND_199 (c6288_wire_301, {c6288_wire_25_15, c6288_wire_117_10});
and_n #(3, 0, 0) AND_200 (c6288_wire_302, {c6288_wire_25_16, c6288_wire_117_11, c6288_wire_303_0});
and_n #(3, 0, 0) AND_201 (c6288_wire_304, {c6288_wire_25_17, c6288_wire_114_11, c6288_wire_305_0});
and_n #(3, 0, 0) AND_202 (c6288_wire_306, {c6288_wire_25_18, c6288_wire_111_11, c6288_wire_307_0});
and_n #(3, 0, 0) AND_203 (c6288_wire_308, {c6288_wire_25_19, c6288_wire_108_11, c6288_wire_309_0});
and_n #(3, 0, 0) AND_204 (c6288_wire_310, {c6288_wire_25_20, c6288_wire_105_11, c6288_wire_311_0});
and_n #(3, 0, 0) AND_205 (c6288_wire_312, {c6288_wire_25_21, c6288_wire_102_11, c6288_wire_313_0});
and_n #(3, 0, 0) AND_206 (c6288_wire_314, {c6288_wire_25_22, c6288_wire_99_11, c6288_wire_315_0});
and_n #(3, 0, 0) AND_207 (c6288_wire_316, {c6288_wire_25_23, c6288_wire_96_11, c6288_wire_317_0});
and_n #(3, 0, 0) AND_208 (c6288_wire_318, {c6288_wire_25_24, c6288_wire_93_11, c6288_wire_319_0});
and_n #(3, 0, 0) AND_209 (c6288_wire_320, {c6288_wire_25_25, c6288_wire_90_11, c6288_wire_321_0});
and_n #(3, 0, 0) AND_210 (c6288_wire_322, {c6288_wire_25_26, c6288_wire_87_11, c6288_wire_323_0});
and_n #(3, 0, 0) AND_211 (c6288_wire_324, {c6288_wire_25_27, c6288_wire_84_11, c6288_wire_325_0});
and_n #(3, 0, 0) AND_212 (c6288_wire_326, {c6288_wire_25_28, c6288_wire_81_11, c6288_wire_327_0});
and_n #(2, 0, 0) AND_213 (c6288_wire_328, {c6288_wire_25_29, c6288_wire_6_28});
and_n #(2, 0, 0) AND_214 (c6288_wire_329, {c6288_wire_330_0, c6288_wire_81_12});
and_n #(2, 0, 0) AND_215 (c6288_wire_331, {c6288_wire_330_1, c6288_wire_84_12});
and_n #(2, 0, 0) AND_216 (c6288_wire_332, {c6288_wire_330_2, c6288_wire_87_12});
and_n #(2, 0, 0) AND_217 (c6288_wire_333, {c6288_wire_330_3, c6288_wire_90_12});
and_n #(2, 0, 0) AND_218 (c6288_wire_334, {c6288_wire_330_4, c6288_wire_93_12});
and_n #(2, 0, 0) AND_219 (c6288_wire_335, {c6288_wire_330_5, c6288_wire_96_12});
and_n #(2, 0, 0) AND_220 (c6288_wire_336, {c6288_wire_330_6, c6288_wire_99_12});
and_n #(2, 0, 0) AND_221 (c6288_wire_337, {c6288_wire_330_7, c6288_wire_102_12});
and_n #(2, 0, 0) AND_222 (c6288_wire_338, {c6288_wire_330_8, c6288_wire_105_12});
and_n #(2, 0, 0) AND_223 (c6288_wire_339, {c6288_wire_330_9, c6288_wire_108_12});
and_n #(2, 0, 0) AND_224 (c6288_wire_340, {c6288_wire_330_10, c6288_wire_111_12});
and_n #(2, 0, 0) AND_225 (c6288_wire_341, {c6288_wire_330_11, c6288_wire_114_12});
and_n #(2, 0, 0) AND_226 (c6288_wire_342, {c6288_wire_330_12, c6288_wire_117_12});
and_n #(2, 0, 0) AND_227 (c6288_wire_343, {c6288_wire_330_13, c6288_wire_114_13});
and_n #(2, 0, 0) AND_228 (c6288_wire_344, {c6288_wire_330_14, c6288_wire_111_13});
and_n #(2, 0, 0) AND_229 (c6288_wire_345, {c6288_wire_330_15, c6288_wire_108_13});
and_n #(2, 0, 0) AND_230 (c6288_wire_346, {c6288_wire_330_16, c6288_wire_105_13});
and_n #(2, 0, 0) AND_231 (c6288_wire_347, {c6288_wire_330_17, c6288_wire_102_13});
and_n #(2, 0, 0) AND_232 (c6288_wire_348, {c6288_wire_330_18, c6288_wire_99_13});
and_n #(2, 0, 0) AND_233 (c6288_wire_349, {c6288_wire_330_19, c6288_wire_96_13});
and_n #(2, 0, 0) AND_234 (c6288_wire_350, {c6288_wire_330_20, c6288_wire_93_13});
and_n #(2, 0, 0) AND_235 (c6288_wire_351, {c6288_wire_330_21, c6288_wire_90_13});
and_n #(2, 0, 0) AND_236 (c6288_wire_352, {c6288_wire_330_22, c6288_wire_87_13});
and_n #(2, 0, 0) AND_237 (c6288_wire_353, {c6288_wire_330_23, c6288_wire_84_13});
and_n #(2, 0, 0) AND_238 (c6288_wire_354, {c6288_wire_330_24, c6288_wire_81_13});
and_n #(2, 0, 0) AND_239 (c6288_wire_355, {c6288_wire_330_25, c6288_wire_6_29});
and_n #(2, 0, 0) AND_240 (c6288_wire_356, {c6288_wire_330_26, c6288_wire_3_15});
and_n #(2, 0, 0) AND_241 (c6288_wire_357, {c6288_wire_330_27, c6288_wire_117_13});
and_n #(2, 0, 0) AND_242 (c6288_wire_358, {c6288_wire_330_28, c6288_wire_359});
and_n #(2, 0, 0) AND_243 (c6288_wire_327, {c6288_wire_330_29, c6288_wire_360});
and_n #(2, 0, 0) AND_244 (c6288_wire_361, {c6288_wire_30_3, c6288_wire_78_12});
and_n #(2, 0, 0) AND_245 (c6288_wire_362, {c6288_wire_30_4, c6288_wire_81_14});
and_n #(2, 0, 0) AND_246 (c6288_wire_363, {c6288_wire_30_5, c6288_wire_84_14});
and_n #(2, 0, 0) AND_247 (c6288_wire_364, {c6288_wire_30_6, c6288_wire_87_14});
and_n #(2, 0, 0) AND_248 (c6288_wire_365, {c6288_wire_30_7, c6288_wire_90_14});
and_n #(2, 0, 0) AND_249 (c6288_wire_366, {c6288_wire_30_8, c6288_wire_93_14});
and_n #(2, 0, 0) AND_250 (c6288_wire_367, {c6288_wire_30_9, c6288_wire_96_14});
and_n #(2, 0, 0) AND_251 (c6288_wire_368, {c6288_wire_30_10, c6288_wire_99_14});
and_n #(2, 0, 0) AND_252 (c6288_wire_369, {c6288_wire_30_11, c6288_wire_102_14});
and_n #(2, 0, 0) AND_253 (c6288_wire_370, {c6288_wire_30_12, c6288_wire_105_14});
and_n #(2, 0, 0) AND_254 (c6288_wire_371, {c6288_wire_30_13, c6288_wire_108_14});
and_n #(2, 0, 0) AND_255 (c6288_wire_372, {c6288_wire_30_14, c6288_wire_111_14});
and_n #(2, 0, 0) AND_256 (c6288_wire_373, {c6288_wire_30_15, c6288_wire_114_14});
and_n #(2, 0, 0) AND_257 (c6288_wire_374, {c6288_wire_30_16, c6288_wire_117_14});
and_n #(3, 0, 0) AND_258 (c6288_wire_375, {c6288_wire_30_17, c6288_wire_117_15, c6288_wire_376_0});
and_n #(3, 0, 0) AND_259 (c6288_wire_377, {c6288_wire_30_18, c6288_wire_114_15, c6288_wire_378_0});
and_n #(3, 0, 0) AND_260 (c6288_wire_379, {c6288_wire_30_19, c6288_wire_111_15, c6288_wire_380_0});
and_n #(3, 0, 0) AND_261 (c6288_wire_381, {c6288_wire_30_20, c6288_wire_108_15, c6288_wire_382_0});
and_n #(3, 0, 0) AND_262 (c6288_wire_383, {c6288_wire_30_21, c6288_wire_105_15, c6288_wire_384_0});
and_n #(3, 0, 0) AND_263 (c6288_wire_385, {c6288_wire_30_22, c6288_wire_102_15, c6288_wire_386_0});
and_n #(3, 0, 0) AND_264 (c6288_wire_387, {c6288_wire_30_23, c6288_wire_99_15, c6288_wire_388_0});
and_n #(3, 0, 0) AND_265 (c6288_wire_389, {c6288_wire_30_24, c6288_wire_96_15, c6288_wire_390_0});
and_n #(3, 0, 0) AND_266 (c6288_wire_391, {c6288_wire_30_25, c6288_wire_93_15, c6288_wire_392_0});
and_n #(3, 0, 0) AND_267 (c6288_wire_393, {c6288_wire_30_26, c6288_wire_90_15, c6288_wire_394_0});
and_n #(3, 0, 0) AND_268 (c6288_wire_395, {c6288_wire_30_27, c6288_wire_87_15, c6288_wire_396_0});
and_n #(3, 0, 0) AND_269 (c6288_wire_397, {c6288_wire_30_28, c6288_wire_84_15, c6288_wire_398_0});
and_n #(3, 0, 0) AND_270 (c6288_wire_399, {c6288_wire_30_29, c6288_wire_81_15, c6288_wire_400_0});
and_n #(3, 0, 0) AND_271 (c6288_wire_401, {c6288_wire_30_30, c6288_wire_78_13, c6288_wire_402_0});
and_n #(2, 0, 0) AND_272 (c6288_wire_403, {c6288_wire_37_3, c6288_wire_78_14});
and_n #(2, 0, 0) AND_273 (c6288_wire_404, {c6288_wire_37_4, c6288_wire_81_16});
and_n #(2, 0, 0) AND_274 (c6288_wire_405, {c6288_wire_37_5, c6288_wire_84_16});
and_n #(2, 0, 0) AND_275 (c6288_wire_406, {c6288_wire_37_6, c6288_wire_87_16});
and_n #(2, 0, 0) AND_276 (c6288_wire_407, {c6288_wire_37_7, c6288_wire_90_16});
and_n #(2, 0, 0) AND_277 (c6288_wire_408, {c6288_wire_37_8, c6288_wire_93_16});
and_n #(2, 0, 0) AND_278 (c6288_wire_409, {c6288_wire_37_9, c6288_wire_96_16});
and_n #(2, 0, 0) AND_279 (c6288_wire_410, {c6288_wire_37_10, c6288_wire_99_16});
and_n #(2, 0, 0) AND_280 (c6288_wire_411, {c6288_wire_37_11, c6288_wire_102_16});
and_n #(2, 0, 0) AND_281 (c6288_wire_412, {c6288_wire_37_12, c6288_wire_105_16});
and_n #(2, 0, 0) AND_282 (c6288_wire_413, {c6288_wire_37_13, c6288_wire_108_16});
and_n #(2, 0, 0) AND_283 (c6288_wire_414, {c6288_wire_37_14, c6288_wire_111_16});
and_n #(2, 0, 0) AND_284 (c6288_wire_415, {c6288_wire_37_15, c6288_wire_114_16});
and_n #(2, 0, 0) AND_285 (c6288_wire_416, {c6288_wire_37_16, c6288_wire_117_16});
and_n #(3, 0, 0) AND_286 (c6288_wire_417, {c6288_wire_37_17, c6288_wire_117_17, c6288_wire_418_0});
and_n #(3, 0, 0) AND_287 (c6288_wire_419, {c6288_wire_37_18, c6288_wire_114_17, c6288_wire_420_0});
and_n #(3, 0, 0) AND_288 (c6288_wire_421, {c6288_wire_37_19, c6288_wire_111_17, c6288_wire_422_0});
and_n #(3, 0, 0) AND_289 (c6288_wire_423, {c6288_wire_37_20, c6288_wire_108_17, c6288_wire_424_0});
and_n #(3, 0, 0) AND_290 (c6288_wire_425, {c6288_wire_37_21, c6288_wire_105_17, c6288_wire_426_0});
and_n #(3, 0, 0) AND_291 (c6288_wire_427, {c6288_wire_37_22, c6288_wire_102_17, c6288_wire_428_0});
and_n #(3, 0, 0) AND_292 (c6288_wire_429, {c6288_wire_37_23, c6288_wire_99_17, c6288_wire_430_0});
and_n #(3, 0, 0) AND_293 (c6288_wire_431, {c6288_wire_37_24, c6288_wire_96_17, c6288_wire_432_0});
and_n #(3, 0, 0) AND_294 (c6288_wire_433, {c6288_wire_37_25, c6288_wire_93_17, c6288_wire_434_0});
and_n #(3, 0, 0) AND_295 (c6288_wire_435, {c6288_wire_37_26, c6288_wire_90_17, c6288_wire_436_0});
and_n #(3, 0, 0) AND_296 (c6288_wire_437, {c6288_wire_37_27, c6288_wire_87_17, c6288_wire_438_0});
and_n #(3, 0, 0) AND_297 (c6288_wire_439, {c6288_wire_37_28, c6288_wire_84_17, c6288_wire_440_0});
and_n #(3, 0, 0) AND_298 (c6288_wire_441, {c6288_wire_37_29, c6288_wire_81_17, c6288_wire_442_0});
and_n #(3, 0, 0) AND_299 (c6288_wire_443, {c6288_wire_37_30, c6288_wire_78_15, c6288_wire_444_0});
and_n #(2, 0, 0) AND_300 (c6288_wire_445, {c6288_wire_42_3, c6288_wire_78_16});
and_n #(2, 0, 0) AND_301 (c6288_wire_446, {c6288_wire_42_4, c6288_wire_81_18});
and_n #(2, 0, 0) AND_302 (c6288_wire_447, {c6288_wire_42_5, c6288_wire_84_18});
and_n #(2, 0, 0) AND_303 (c6288_wire_448, {c6288_wire_42_6, c6288_wire_87_18});
and_n #(2, 0, 0) AND_304 (c6288_wire_449, {c6288_wire_42_7, c6288_wire_90_18});
and_n #(2, 0, 0) AND_305 (c6288_wire_450, {c6288_wire_42_8, c6288_wire_93_18});
and_n #(2, 0, 0) AND_306 (c6288_wire_451, {c6288_wire_42_9, c6288_wire_96_18});
and_n #(2, 0, 0) AND_307 (c6288_wire_452, {c6288_wire_42_10, c6288_wire_99_18});
and_n #(2, 0, 0) AND_308 (c6288_wire_453, {c6288_wire_42_11, c6288_wire_102_18});
and_n #(2, 0, 0) AND_309 (c6288_wire_454, {c6288_wire_42_12, c6288_wire_105_18});
and_n #(2, 0, 0) AND_310 (c6288_wire_455, {c6288_wire_42_13, c6288_wire_108_18});
and_n #(2, 0, 0) AND_311 (c6288_wire_456, {c6288_wire_42_14, c6288_wire_111_18});
and_n #(2, 0, 0) AND_312 (c6288_wire_457, {c6288_wire_42_15, c6288_wire_114_18});
and_n #(2, 0, 0) AND_313 (c6288_wire_458, {c6288_wire_42_16, c6288_wire_117_18});
and_n #(3, 0, 0) AND_314 (c6288_wire_459, {c6288_wire_42_17, c6288_wire_117_19, c6288_wire_460_0});
and_n #(3, 0, 0) AND_315 (c6288_wire_461, {c6288_wire_42_18, c6288_wire_114_19, c6288_wire_462_0});
and_n #(3, 0, 0) AND_316 (c6288_wire_463, {c6288_wire_42_19, c6288_wire_111_19, c6288_wire_464_0});
and_n #(3, 0, 0) AND_317 (c6288_wire_465, {c6288_wire_42_20, c6288_wire_108_19, c6288_wire_466_0});
and_n #(3, 0, 0) AND_318 (c6288_wire_467, {c6288_wire_42_21, c6288_wire_105_19, c6288_wire_468_0});
and_n #(3, 0, 0) AND_319 (c6288_wire_469, {c6288_wire_42_22, c6288_wire_102_19, c6288_wire_470_0});
and_n #(3, 0, 0) AND_320 (c6288_wire_471, {c6288_wire_42_23, c6288_wire_99_19, c6288_wire_472_0});
and_n #(3, 0, 0) AND_321 (c6288_wire_473, {c6288_wire_42_24, c6288_wire_96_19, c6288_wire_474_0});
and_n #(3, 0, 0) AND_322 (c6288_wire_475, {c6288_wire_42_25, c6288_wire_93_19, c6288_wire_476_0});
and_n #(3, 0, 0) AND_323 (c6288_wire_477, {c6288_wire_42_26, c6288_wire_90_19, c6288_wire_478_0});
and_n #(3, 0, 0) AND_324 (c6288_wire_479, {c6288_wire_42_27, c6288_wire_87_19, c6288_wire_480_0});
and_n #(3, 0, 0) AND_325 (c6288_wire_481, {c6288_wire_42_28, c6288_wire_84_19, c6288_wire_482_0});
and_n #(3, 0, 0) AND_326 (c6288_wire_483, {c6288_wire_42_29, c6288_wire_81_19, c6288_wire_484_0});
and_n #(3, 0, 0) AND_327 (c6288_wire_485, {c6288_wire_42_30, c6288_wire_78_17, c6288_wire_486_0});
and_n #(2, 0, 0) AND_328 (c6288_wire_487, {c6288_wire_47_3, c6288_wire_78_18});
and_n #(2, 0, 0) AND_329 (c6288_wire_488, {c6288_wire_47_4, c6288_wire_81_20});
and_n #(2, 0, 0) AND_330 (c6288_wire_489, {c6288_wire_47_5, c6288_wire_84_20});
and_n #(2, 0, 0) AND_331 (c6288_wire_490, {c6288_wire_47_6, c6288_wire_87_20});
and_n #(2, 0, 0) AND_332 (c6288_wire_491, {c6288_wire_47_7, c6288_wire_90_20});
and_n #(2, 0, 0) AND_333 (c6288_wire_492, {c6288_wire_47_8, c6288_wire_93_20});
and_n #(2, 0, 0) AND_334 (c6288_wire_493, {c6288_wire_47_9, c6288_wire_96_20});
and_n #(2, 0, 0) AND_335 (c6288_wire_494, {c6288_wire_47_10, c6288_wire_99_20});
and_n #(2, 0, 0) AND_336 (c6288_wire_495, {c6288_wire_47_11, c6288_wire_102_20});
and_n #(2, 0, 0) AND_337 (c6288_wire_496, {c6288_wire_47_12, c6288_wire_105_20});
and_n #(2, 0, 0) AND_338 (c6288_wire_497, {c6288_wire_47_13, c6288_wire_108_20});
and_n #(2, 0, 0) AND_339 (c6288_wire_498, {c6288_wire_47_14, c6288_wire_111_20});
and_n #(2, 0, 0) AND_340 (c6288_wire_499, {c6288_wire_47_15, c6288_wire_114_20});
and_n #(2, 0, 0) AND_341 (c6288_wire_500, {c6288_wire_47_16, c6288_wire_117_20});
and_n #(3, 0, 0) AND_342 (c6288_wire_501, {c6288_wire_47_17, c6288_wire_117_21, c6288_wire_502_0});
and_n #(3, 0, 0) AND_343 (c6288_wire_503, {c6288_wire_47_18, c6288_wire_114_21, c6288_wire_504_0});
and_n #(3, 0, 0) AND_344 (c6288_wire_505, {c6288_wire_47_19, c6288_wire_111_21, c6288_wire_506_0});
and_n #(3, 0, 0) AND_345 (c6288_wire_507, {c6288_wire_47_20, c6288_wire_108_21, c6288_wire_508_0});
and_n #(3, 0, 0) AND_346 (c6288_wire_509, {c6288_wire_47_21, c6288_wire_105_21, c6288_wire_510_0});
and_n #(3, 0, 0) AND_347 (c6288_wire_511, {c6288_wire_47_22, c6288_wire_102_21, c6288_wire_512_0});
and_n #(3, 0, 0) AND_348 (c6288_wire_513, {c6288_wire_47_23, c6288_wire_99_21, c6288_wire_514_0});
and_n #(3, 0, 0) AND_349 (c6288_wire_515, {c6288_wire_47_24, c6288_wire_96_21, c6288_wire_516_0});
and_n #(3, 0, 0) AND_350 (c6288_wire_517, {c6288_wire_47_25, c6288_wire_93_21, c6288_wire_518_0});
and_n #(3, 0, 0) AND_351 (c6288_wire_519, {c6288_wire_47_26, c6288_wire_90_21, c6288_wire_520_0});
and_n #(3, 0, 0) AND_352 (c6288_wire_521, {c6288_wire_47_27, c6288_wire_87_21, c6288_wire_522_0});
and_n #(3, 0, 0) AND_353 (c6288_wire_523, {c6288_wire_47_28, c6288_wire_84_21, c6288_wire_524_0});
and_n #(3, 0, 0) AND_354 (c6288_wire_525, {c6288_wire_47_29, c6288_wire_81_21, c6288_wire_526_0});
and_n #(3, 0, 0) AND_355 (c6288_wire_527, {c6288_wire_47_30, c6288_wire_78_19, c6288_wire_528_0});
and_n #(2, 0, 0) AND_356 (c6288_wire_529, {c6288_wire_52_3, c6288_wire_78_20});
and_n #(2, 0, 0) AND_357 (c6288_wire_530, {c6288_wire_52_4, c6288_wire_81_22});
and_n #(2, 0, 0) AND_358 (c6288_wire_531, {c6288_wire_52_5, c6288_wire_84_22});
and_n #(2, 0, 0) AND_359 (c6288_wire_532, {c6288_wire_52_6, c6288_wire_87_22});
and_n #(2, 0, 0) AND_360 (c6288_wire_533, {c6288_wire_52_7, c6288_wire_90_22});
and_n #(2, 0, 0) AND_361 (c6288_wire_534, {c6288_wire_52_8, c6288_wire_93_22});
and_n #(2, 0, 0) AND_362 (c6288_wire_535, {c6288_wire_52_9, c6288_wire_96_22});
and_n #(2, 0, 0) AND_363 (c6288_wire_536, {c6288_wire_52_10, c6288_wire_99_22});
and_n #(2, 0, 0) AND_364 (c6288_wire_537, {c6288_wire_52_11, c6288_wire_102_22});
and_n #(2, 0, 0) AND_365 (c6288_wire_538, {c6288_wire_52_12, c6288_wire_105_22});
and_n #(2, 0, 0) AND_366 (c6288_wire_539, {c6288_wire_52_13, c6288_wire_108_22});
and_n #(2, 0, 0) AND_367 (c6288_wire_540, {c6288_wire_52_14, c6288_wire_111_22});
and_n #(2, 0, 0) AND_368 (c6288_wire_541, {c6288_wire_52_15, c6288_wire_114_22});
and_n #(2, 0, 0) AND_369 (c6288_wire_542, {c6288_wire_52_16, c6288_wire_117_22});
and_n #(3, 0, 0) AND_370 (c6288_wire_543, {c6288_wire_52_17, c6288_wire_117_23, c6288_wire_544_0});
and_n #(3, 0, 0) AND_371 (c6288_wire_545, {c6288_wire_52_18, c6288_wire_114_23, c6288_wire_546_0});
and_n #(3, 0, 0) AND_372 (c6288_wire_547, {c6288_wire_52_19, c6288_wire_111_23, c6288_wire_548_0});
and_n #(3, 0, 0) AND_373 (c6288_wire_549, {c6288_wire_52_20, c6288_wire_108_23, c6288_wire_550_0});
and_n #(3, 0, 0) AND_374 (c6288_wire_551, {c6288_wire_52_21, c6288_wire_105_23, c6288_wire_552_0});
and_n #(3, 0, 0) AND_375 (c6288_wire_553, {c6288_wire_52_22, c6288_wire_102_23, c6288_wire_554_0});
and_n #(3, 0, 0) AND_376 (c6288_wire_555, {c6288_wire_52_23, c6288_wire_99_23, c6288_wire_556_0});
and_n #(3, 0, 0) AND_377 (c6288_wire_557, {c6288_wire_52_24, c6288_wire_96_23, c6288_wire_558_0});
and_n #(3, 0, 0) AND_378 (c6288_wire_559, {c6288_wire_52_25, c6288_wire_93_23, c6288_wire_560_0});
and_n #(3, 0, 0) AND_379 (c6288_wire_561, {c6288_wire_52_26, c6288_wire_90_23, c6288_wire_562_0});
and_n #(3, 0, 0) AND_380 (c6288_wire_563, {c6288_wire_52_27, c6288_wire_87_23, c6288_wire_564_0});
and_n #(3, 0, 0) AND_381 (c6288_wire_565, {c6288_wire_52_28, c6288_wire_84_23, c6288_wire_566_0});
and_n #(3, 0, 0) AND_382 (c6288_wire_567, {c6288_wire_52_29, c6288_wire_81_23, c6288_wire_568_0});
and_n #(3, 0, 0) AND_383 (c6288_wire_569, {c6288_wire_52_30, c6288_wire_78_21, c6288_wire_570_0});
and_n #(2, 0, 0) AND_384 (c6288_wire_571, {c6288_wire_57_3, c6288_wire_78_22});
and_n #(2, 0, 0) AND_385 (c6288_wire_572, {c6288_wire_57_4, c6288_wire_81_24});
and_n #(2, 0, 0) AND_386 (c6288_wire_573, {c6288_wire_57_5, c6288_wire_84_24});
and_n #(2, 0, 0) AND_387 (c6288_wire_574, {c6288_wire_57_6, c6288_wire_87_24});
and_n #(2, 0, 0) AND_388 (c6288_wire_575, {c6288_wire_57_7, c6288_wire_90_24});
and_n #(2, 0, 0) AND_389 (c6288_wire_576, {c6288_wire_57_8, c6288_wire_93_24});
and_n #(2, 0, 0) AND_390 (c6288_wire_577, {c6288_wire_57_9, c6288_wire_96_24});
and_n #(2, 0, 0) AND_391 (c6288_wire_578, {c6288_wire_57_10, c6288_wire_99_24});
and_n #(2, 0, 0) AND_392 (c6288_wire_579, {c6288_wire_57_11, c6288_wire_102_24});
and_n #(2, 0, 0) AND_393 (c6288_wire_580, {c6288_wire_57_12, c6288_wire_105_24});
and_n #(2, 0, 0) AND_394 (c6288_wire_581, {c6288_wire_57_13, c6288_wire_108_24});
and_n #(2, 0, 0) AND_395 (c6288_wire_582, {c6288_wire_57_14, c6288_wire_111_24});
and_n #(2, 0, 0) AND_396 (c6288_wire_583, {c6288_wire_57_15, c6288_wire_114_24});
and_n #(2, 0, 0) AND_397 (c6288_wire_584, {c6288_wire_57_16, c6288_wire_117_24});
and_n #(3, 0, 0) AND_398 (c6288_wire_585, {c6288_wire_57_17, c6288_wire_117_25, c6288_wire_586_0});
and_n #(3, 0, 0) AND_399 (c6288_wire_587, {c6288_wire_57_18, c6288_wire_114_25, c6288_wire_588_0});
and_n #(3, 0, 0) AND_400 (c6288_wire_589, {c6288_wire_57_19, c6288_wire_111_25, c6288_wire_590_0});
and_n #(3, 0, 0) AND_401 (c6288_wire_591, {c6288_wire_57_20, c6288_wire_108_25, c6288_wire_592_0});
and_n #(3, 0, 0) AND_402 (c6288_wire_593, {c6288_wire_57_21, c6288_wire_105_25, c6288_wire_594_0});
and_n #(3, 0, 0) AND_403 (c6288_wire_595, {c6288_wire_57_22, c6288_wire_102_25, c6288_wire_596_0});
and_n #(3, 0, 0) AND_404 (c6288_wire_597, {c6288_wire_57_23, c6288_wire_99_25, c6288_wire_598_0});
and_n #(3, 0, 0) AND_405 (c6288_wire_599, {c6288_wire_57_24, c6288_wire_96_25, c6288_wire_600_0});
and_n #(3, 0, 0) AND_406 (c6288_wire_601, {c6288_wire_57_25, c6288_wire_93_25, c6288_wire_602_0});
and_n #(3, 0, 0) AND_407 (c6288_wire_603, {c6288_wire_57_26, c6288_wire_90_25, c6288_wire_604_0});
and_n #(3, 0, 0) AND_408 (c6288_wire_605, {c6288_wire_57_27, c6288_wire_87_25, c6288_wire_606_0});
and_n #(3, 0, 0) AND_409 (c6288_wire_607, {c6288_wire_57_28, c6288_wire_84_25, c6288_wire_608_0});
and_n #(3, 0, 0) AND_410 (c6288_wire_609, {c6288_wire_57_29, c6288_wire_81_25, c6288_wire_610_0});
and_n #(3, 0, 0) AND_411 (c6288_wire_611, {c6288_wire_57_30, c6288_wire_78_23, c6288_wire_612_0});
and_n #(2, 0, 0) AND_412 (c6288_wire_613, {c6288_wire_62_3, c6288_wire_78_24});
and_n #(2, 0, 0) AND_413 (c6288_wire_614, {c6288_wire_62_4, c6288_wire_81_26});
and_n #(2, 0, 0) AND_414 (c6288_wire_615, {c6288_wire_62_5, c6288_wire_84_26});
and_n #(2, 0, 0) AND_415 (c6288_wire_616, {c6288_wire_62_6, c6288_wire_87_26});
and_n #(2, 0, 0) AND_416 (c6288_wire_617, {c6288_wire_62_7, c6288_wire_90_26});
and_n #(2, 0, 0) AND_417 (c6288_wire_618, {c6288_wire_62_8, c6288_wire_93_26});
and_n #(2, 0, 0) AND_418 (c6288_wire_619, {c6288_wire_62_9, c6288_wire_96_26});
and_n #(2, 0, 0) AND_419 (c6288_wire_620, {c6288_wire_62_10, c6288_wire_99_26});
and_n #(2, 0, 0) AND_420 (c6288_wire_621, {c6288_wire_62_11, c6288_wire_102_26});
and_n #(2, 0, 0) AND_421 (c6288_wire_622, {c6288_wire_62_12, c6288_wire_105_26});
and_n #(2, 0, 0) AND_422 (c6288_wire_623, {c6288_wire_62_13, c6288_wire_108_26});
and_n #(2, 0, 0) AND_423 (c6288_wire_624, {c6288_wire_62_14, c6288_wire_111_26});
and_n #(2, 0, 0) AND_424 (c6288_wire_625, {c6288_wire_62_15, c6288_wire_114_26});
and_n #(2, 0, 0) AND_425 (c6288_wire_626, {c6288_wire_62_16, c6288_wire_117_26});
and_n #(3, 0, 0) AND_426 (c6288_wire_627, {c6288_wire_62_17, c6288_wire_117_27, c6288_wire_628_0});
and_n #(3, 0, 0) AND_427 (c6288_wire_629, {c6288_wire_62_18, c6288_wire_114_27, c6288_wire_630_0});
and_n #(3, 0, 0) AND_428 (c6288_wire_631, {c6288_wire_62_19, c6288_wire_111_27, c6288_wire_632_0});
and_n #(3, 0, 0) AND_429 (c6288_wire_633, {c6288_wire_62_20, c6288_wire_108_27, c6288_wire_634_0});
and_n #(3, 0, 0) AND_430 (c6288_wire_635, {c6288_wire_62_21, c6288_wire_105_27, c6288_wire_636_0});
and_n #(3, 0, 0) AND_431 (c6288_wire_637, {c6288_wire_62_22, c6288_wire_102_27, c6288_wire_638_0});
and_n #(3, 0, 0) AND_432 (c6288_wire_639, {c6288_wire_62_23, c6288_wire_99_27, c6288_wire_640_0});
and_n #(3, 0, 0) AND_433 (c6288_wire_641, {c6288_wire_62_24, c6288_wire_96_27, c6288_wire_642_0});
and_n #(3, 0, 0) AND_434 (c6288_wire_643, {c6288_wire_62_25, c6288_wire_93_27, c6288_wire_644_0});
and_n #(3, 0, 0) AND_435 (c6288_wire_645, {c6288_wire_62_26, c6288_wire_90_27, c6288_wire_646_0});
and_n #(3, 0, 0) AND_436 (c6288_wire_647, {c6288_wire_62_27, c6288_wire_87_27, c6288_wire_648_0});
and_n #(3, 0, 0) AND_437 (c6288_wire_649, {c6288_wire_62_28, c6288_wire_84_27, c6288_wire_650_0});
and_n #(3, 0, 0) AND_438 (c6288_wire_651, {c6288_wire_62_29, c6288_wire_81_27, c6288_wire_652_0});
and_n #(3, 0, 0) AND_439 (c6288_wire_653, {c6288_wire_62_30, c6288_wire_78_25, c6288_wire_654_0});
and_n #(2, 0, 0) AND_440 (c6288_wire_655, {c6288_wire_67_3, c6288_wire_78_26});
and_n #(2, 0, 0) AND_441 (c6288_wire_656, {c6288_wire_67_4, c6288_wire_81_28});
and_n #(2, 0, 0) AND_442 (c6288_wire_657, {c6288_wire_67_5, c6288_wire_84_28});
and_n #(2, 0, 0) AND_443 (c6288_wire_658, {c6288_wire_67_6, c6288_wire_87_28});
and_n #(2, 0, 0) AND_444 (c6288_wire_659, {c6288_wire_67_7, c6288_wire_90_28});
and_n #(2, 0, 0) AND_445 (c6288_wire_660, {c6288_wire_67_8, c6288_wire_93_28});
and_n #(2, 0, 0) AND_446 (c6288_wire_661, {c6288_wire_67_9, c6288_wire_96_28});
and_n #(2, 0, 0) AND_447 (c6288_wire_662, {c6288_wire_67_10, c6288_wire_99_28});
and_n #(2, 0, 0) AND_448 (c6288_wire_663, {c6288_wire_67_11, c6288_wire_102_28});
and_n #(2, 0, 0) AND_449 (c6288_wire_664, {c6288_wire_67_12, c6288_wire_105_28});
and_n #(2, 0, 0) AND_450 (c6288_wire_665, {c6288_wire_67_13, c6288_wire_108_28});
and_n #(2, 0, 0) AND_451 (c6288_wire_666, {c6288_wire_67_14, c6288_wire_111_28});
and_n #(2, 0, 0) AND_452 (c6288_wire_667, {c6288_wire_67_15, c6288_wire_114_28});
and_n #(2, 0, 0) AND_453 (c6288_wire_668, {c6288_wire_67_16, c6288_wire_117_28});
and_n #(3, 0, 0) AND_454 (c6288_wire_669, {c6288_wire_67_17, c6288_wire_117_29, c6288_wire_670_0});
and_n #(3, 0, 0) AND_455 (c6288_wire_671, {c6288_wire_67_18, c6288_wire_114_29, c6288_wire_672_0});
and_n #(3, 0, 0) AND_456 (c6288_wire_673, {c6288_wire_67_19, c6288_wire_111_29, c6288_wire_674_0});
and_n #(3, 0, 0) AND_457 (c6288_wire_675, {c6288_wire_67_20, c6288_wire_108_29, c6288_wire_676_0});
and_n #(3, 0, 0) AND_458 (c6288_wire_677, {c6288_wire_67_21, c6288_wire_105_29, c6288_wire_678_0});
and_n #(3, 0, 0) AND_459 (c6288_wire_679, {c6288_wire_67_22, c6288_wire_102_29, c6288_wire_680_0});
and_n #(3, 0, 0) AND_460 (c6288_wire_681, {c6288_wire_67_23, c6288_wire_99_29, c6288_wire_682_0});
and_n #(3, 0, 0) AND_461 (c6288_wire_683, {c6288_wire_67_24, c6288_wire_96_29, c6288_wire_684_0});
and_n #(3, 0, 0) AND_462 (c6288_wire_685, {c6288_wire_67_25, c6288_wire_93_29, c6288_wire_686_0});
and_n #(3, 0, 0) AND_463 (c6288_wire_687, {c6288_wire_67_26, c6288_wire_90_29, c6288_wire_688_0});
and_n #(3, 0, 0) AND_464 (c6288_wire_689, {c6288_wire_67_27, c6288_wire_87_29, c6288_wire_690_0});
and_n #(3, 0, 0) AND_465 (c6288_wire_691, {c6288_wire_67_28, c6288_wire_84_29, c6288_wire_692_0});
and_n #(3, 0, 0) AND_466 (c6288_wire_693, {c6288_wire_67_29, c6288_wire_81_29, c6288_wire_694_0});
and_n #(3, 0, 0) AND_467 (c6288_wire_695, {c6288_wire_67_30, c6288_wire_78_27, c6288_wire_696_0});
and_n #(2, 0, 0) AND_468 (c6288_wire_697, {c6288_wire_5_3, c6288_wire_78_28});
and_n #(2, 0, 0) AND_469 (c6288_wire_698, {c6288_wire_5_4, c6288_wire_81_30});
and_n #(2, 0, 0) AND_470 (c6288_wire_699, {c6288_wire_5_5, c6288_wire_84_30});
and_n #(2, 0, 0) AND_471 (c6288_wire_700, {c6288_wire_5_6, c6288_wire_87_30});
and_n #(2, 0, 0) AND_472 (c6288_wire_701, {c6288_wire_5_7, c6288_wire_90_30});
and_n #(2, 0, 0) AND_473 (c6288_wire_702, {c6288_wire_5_8, c6288_wire_93_30});
and_n #(2, 0, 0) AND_474 (c6288_wire_703, {c6288_wire_5_9, c6288_wire_96_30});
and_n #(2, 0, 0) AND_475 (c6288_wire_704, {c6288_wire_5_10, c6288_wire_99_30});
and_n #(2, 0, 0) AND_476 (c6288_wire_705, {c6288_wire_5_11, c6288_wire_102_30});
and_n #(2, 0, 0) AND_477 (c6288_wire_706, {c6288_wire_5_12, c6288_wire_105_30});
and_n #(2, 0, 0) AND_478 (c6288_wire_707, {c6288_wire_5_13, c6288_wire_108_30});
and_n #(2, 0, 0) AND_479 (c6288_wire_708, {c6288_wire_5_14, c6288_wire_111_30});
and_n #(2, 0, 0) AND_480 (c6288_wire_709, {c6288_wire_5_15, c6288_wire_114_30});
and_n #(2, 0, 0) AND_481 (c6288_wire_710, {c6288_wire_5_16, c6288_wire_117_30});
and_n #(3, 0, 0) AND_482 (c6288_wire_711, {c6288_wire_5_17, c6288_wire_117_31, c6288_wire_712_0});
and_n #(3, 0, 0) AND_483 (c6288_wire_713, {c6288_wire_5_18, c6288_wire_114_31, c6288_wire_714_0});
and_n #(3, 0, 0) AND_484 (c6288_wire_715, {c6288_wire_5_19, c6288_wire_111_31, c6288_wire_716_0});
and_n #(3, 0, 0) AND_485 (c6288_wire_717, {c6288_wire_5_20, c6288_wire_108_31, c6288_wire_718_0});
and_n #(3, 0, 0) AND_486 (c6288_wire_719, {c6288_wire_5_21, c6288_wire_105_31, c6288_wire_720_0});
and_n #(3, 0, 0) AND_487 (c6288_wire_721, {c6288_wire_5_22, c6288_wire_102_31, c6288_wire_722_0});
and_n #(3, 0, 0) AND_488 (c6288_wire_723, {c6288_wire_5_23, c6288_wire_99_31, c6288_wire_724_0});
and_n #(3, 0, 0) AND_489 (c6288_wire_725, {c6288_wire_5_24, c6288_wire_96_31, c6288_wire_726_0});
and_n #(3, 0, 0) AND_490 (c6288_wire_727, {c6288_wire_5_25, c6288_wire_93_31, c6288_wire_728_0});
and_n #(3, 0, 0) AND_491 (c6288_wire_729, {c6288_wire_5_26, c6288_wire_90_31, c6288_wire_730_0});
and_n #(3, 0, 0) AND_492 (c6288_wire_731, {c6288_wire_5_27, c6288_wire_87_31, c6288_wire_732_0});
and_n #(3, 0, 0) AND_493 (c6288_wire_733, {c6288_wire_5_28, c6288_wire_84_31, c6288_wire_734_0});
and_n #(3, 0, 0) AND_494 (c6288_wire_735, {c6288_wire_5_29, c6288_wire_81_31, c6288_wire_736_0});
and_n #(3, 0, 0) AND_495 (c6288_wire_737, {c6288_wire_5_30, c6288_wire_78_29, c6288_wire_738_0});
and_n #(2, 0, 0) AND_496 (c6288_wire_739, {c6288_wire_6_30, c6288_wire_740_0});
and_n #(2, 0, 0) AND_497 (c6288_wire_741, {c6288_wire_6_31, c6288_wire_740_1});
or_n #(2, 0, 0) OR_1 (c6288_wire_359, {c6288_wire_78_30, c6288_wire_739});
notg #(0, 0) NOT_15 (c6288_wire_742, c6288_wire_78_31);
and_n #(2, 0, 0) AND_498 (c6288_wire_743, {c6288_wire_78_32, c6288_wire_744});
and_n #(2, 0, 0) AND_499 (c6288_wire_745, {c6288_wire_31_0, c6288_wire_746_0});
notg #(0, 0) NOT_16 (c6288_wire_747, c6288_wire_31_1);
xor_n #(2, 0, 0) XOR_1 (c6288_wire_748, {c6288_wire_749_0, c6288_wire_750_0});
or_n #(2, 0, 0) OR_2 (c6288_wire_749, {c6288_wire_751, c6288_wire_752});
and_n #(2, 0, 0) AND_500 (c6288_wire_753, {c6288_wire_749_1, c6288_wire_750_1});
and_n #(2, 0, 0) AND_501 (c6288_wire_751, {c6288_wire_754_0, c6288_wire_755_0});
notg #(0, 0) NOT_17 (c6288_wire_752, c6288_wire_756_0);
xor_n #(2, 0, 0) XOR_2 (c6288_wire_757, {c6288_wire_758_0, c6288_wire_759_0});
or_n #(2, 0, 0) OR_3 (c6288_wire_758, {c6288_wire_753, c6288_wire_760});
and_n #(2, 0, 0) AND_502 (c6288_wire_761, {c6288_wire_758_1, c6288_wire_759_1});
notg #(0, 0) NOT_18 (c6288_wire_760, c6288_wire_762_0);
xor_n #(2, 0, 0) XOR_3 (c6288_wire_763, {c6288_wire_764_0, c6288_wire_765_0});
or_n #(2, 0, 0) OR_4 (c6288_wire_764, {c6288_wire_761, c6288_wire_766});
and_n #(2, 0, 0) AND_503 (c6288_wire_767, {c6288_wire_764_1, c6288_wire_765_1});
notg #(0, 0) NOT_19 (c6288_wire_766, c6288_wire_768_0);
xor_n #(2, 0, 0) XOR_4 (c6288_wire_769, {c6288_wire_770_0, c6288_wire_771_0});
or_n #(2, 0, 0) OR_5 (c6288_wire_770, {c6288_wire_767, c6288_wire_772});
and_n #(2, 0, 0) AND_504 (c6288_wire_773, {c6288_wire_770_1, c6288_wire_771_1});
notg #(0, 0) NOT_20 (c6288_wire_772, c6288_wire_774_0);
xor_n #(2, 0, 0) XOR_5 (c6288_wire_775, {c6288_wire_776_0, c6288_wire_777_0});
or_n #(2, 0, 0) OR_6 (c6288_wire_776, {c6288_wire_773, c6288_wire_778});
notg #(0, 0) NOT_21 (c6288_wire_778, c6288_wire_779_0);
nor_n #(2, 0, 0) NOR_1 (c6288_wire_780, {c6288_wire_776_1, c6288_wire_777_1});
xor_n #(2, 0, 0) XOR_6 (c6288_wire_781, {c6288_wire_780_0, c6288_wire_782_0});
notg #(0, 0) NOT_22 (c6288_wire_783, c6288_wire_780_1);
xor_n #(2, 0, 0) XOR_7 (c6288_wire_784, {c6288_wire_785_0, c6288_wire_786_0});
or_n #(2, 0, 0) OR_7 (c6288_wire_785, {c6288_wire_787, c6288_wire_788});
and_n #(2, 0, 0) AND_505 (c6288_wire_789, {c6288_wire_785_1, c6288_wire_786_1});
and_n #(2, 0, 0) AND_506 (c6288_wire_788, {c6288_wire_747, c6288_wire_746_1});
notg #(0, 0) NOT_23 (c6288_wire_787, c6288_wire_790_0);
xor_n #(2, 0, 0) XOR_8 (c6288_wire_791, {c6288_wire_792_0, c6288_wire_793_0});
or_n #(2, 0, 0) OR_8 (c6288_wire_792, {c6288_wire_789, c6288_wire_794});
and_n #(2, 0, 0) AND_507 (c6288_wire_795, {c6288_wire_792_1, c6288_wire_793_1});
notg #(0, 0) NOT_24 (c6288_wire_794, c6288_wire_796_0);
xor_n #(2, 0, 0) XOR_9 (c6288_wire_797, {c6288_wire_798_0, c6288_wire_799_0});
or_n #(2, 0, 0) OR_9 (c6288_wire_798, {c6288_wire_795, c6288_wire_800});
and_n #(2, 0, 0) AND_508 (c6288_wire_801, {c6288_wire_798_1, c6288_wire_799_1});
notg #(0, 0) NOT_25 (c6288_wire_800, c6288_wire_802_0);
xor_n #(2, 0, 0) XOR_10 (c6288_wire_803, {c6288_wire_804_0, c6288_wire_805_0});
or_n #(2, 0, 0) OR_10 (c6288_wire_804, {c6288_wire_801, c6288_wire_806});
and_n #(2, 0, 0) AND_509 (c6288_wire_807, {c6288_wire_804_1, c6288_wire_805_1});
notg #(0, 0) NOT_26 (c6288_wire_806, c6288_wire_808_0);
xor_n #(2, 0, 0) XOR_11 (c6288_wire_809, {c6288_wire_810_0, c6288_wire_811_0});
or_n #(2, 0, 0) OR_11 (c6288_wire_810, {c6288_wire_807, c6288_wire_812});
and_n #(2, 0, 0) AND_510 (c6288_wire_813, {c6288_wire_810_1, c6288_wire_811_1});
notg #(0, 0) NOT_27 (c6288_wire_812, c6288_wire_814_0);
xor_n #(2, 0, 0) XOR_12 (c6288_wire_815, {c6288_wire_816_0, c6288_wire_817_0});
or_n #(2, 0, 0) OR_12 (c6288_wire_816, {c6288_wire_813, c6288_wire_818});
and_n #(2, 0, 0) AND_511 (c6288_wire_819, {c6288_wire_816_1, c6288_wire_817_1});
notg #(0, 0) NOT_28 (c6288_wire_818, c6288_wire_820_0);
xor_n #(2, 0, 0) XOR_13 (c6288_wire_821, {c6288_wire_822_0, c6288_wire_823_0});
or_n #(2, 0, 0) OR_13 (c6288_wire_822, {c6288_wire_819, c6288_wire_824});
and_n #(2, 0, 0) AND_512 (c6288_wire_825, {c6288_wire_822_1, c6288_wire_823_1});
notg #(0, 0) NOT_29 (c6288_wire_824, c6288_wire_826_0);
xor_n #(2, 0, 0) XOR_14 (c6288_wire_827, {c6288_wire_828_0, c6288_wire_829_0});
or_n #(2, 0, 0) OR_14 (c6288_wire_828, {c6288_wire_825, c6288_wire_830});
and_n #(2, 0, 0) AND_513 (c6288_wire_831, {c6288_wire_828_1, c6288_wire_829_1});
notg #(0, 0) NOT_30 (c6288_wire_830, c6288_wire_832_0);
xor_n #(2, 0, 0) XOR_15 (c6288_wire_833, {c6288_wire_754_1, c6288_wire_755_1});
or_n #(2, 0, 0) OR_15 (c6288_wire_754, {c6288_wire_831, c6288_wire_834});
notg #(0, 0) NOT_31 (c6288_wire_834, c6288_wire_835_0);
and_n #(2, 0, 0) AND_514 (c6288_wire_836, {c6288_wire_11_0, c6288_wire_837_0});
notg #(0, 0) NOT_32 (c6288_wire_838, c6288_wire_11_1);
xor_n #(2, 0, 0) XOR_16 (c6288_wire_140, {c6288_wire_839_0, c6288_wire_840_0});
or_n #(2, 0, 0) OR_16 (c6288_wire_839, {c6288_wire_841, c6288_wire_842});
and_n #(2, 0, 0) AND_515 (c6288_wire_843, {c6288_wire_839_1, c6288_wire_840_1});
and_n #(2, 0, 0) AND_516 (c6288_wire_841, {c6288_wire_844_0, c6288_wire_845_0});
notg #(0, 0) NOT_33 (c6288_wire_842, c6288_wire_846);
xor_n #(2, 0, 0) XOR_17 (c6288_wire_138, {c6288_wire_847_0, c6288_wire_848_0});
or_n #(2, 0, 0) OR_17 (c6288_wire_847, {c6288_wire_843, c6288_wire_849});
and_n #(2, 0, 0) AND_517 (c6288_wire_850, {c6288_wire_847_1, c6288_wire_848_1});
notg #(0, 0) NOT_34 (c6288_wire_849, c6288_wire_851);
xor_n #(2, 0, 0) XOR_18 (c6288_wire_136, {c6288_wire_852_0, c6288_wire_853_0});
or_n #(2, 0, 0) OR_18 (c6288_wire_852, {c6288_wire_850, c6288_wire_854});
and_n #(2, 0, 0) AND_518 (c6288_wire_855, {c6288_wire_852_1, c6288_wire_853_1});
notg #(0, 0) NOT_35 (c6288_wire_854, c6288_wire_856);
xor_n #(2, 0, 0) XOR_19 (c6288_wire_134, {c6288_wire_857_0, c6288_wire_858_0});
or_n #(2, 0, 0) OR_19 (c6288_wire_857, {c6288_wire_855, c6288_wire_859});
and_n #(2, 0, 0) AND_519 (c6288_wire_860, {c6288_wire_857_1, c6288_wire_858_1});
notg #(0, 0) NOT_36 (c6288_wire_859, c6288_wire_861);
xor_n #(2, 0, 0) XOR_20 (c6288_wire_862, {c6288_wire_863_0, c6288_wire_864_0});
or_n #(2, 0, 0) OR_20 (c6288_wire_863, {c6288_wire_860, c6288_wire_865});
and_n #(2, 0, 0) AND_520 (c6288_wire_866, {c6288_wire_863_1, c6288_wire_864_1});
notg #(0, 0) NOT_37 (c6288_wire_865, c6288_wire_867);
and_n #(2, 0, 0) AND_521 (c6288_wire_868, {c6288_wire_869_0, c6288_wire_870_0});
or_n #(2, 0, 0) OR_21 (c6288_wire_869, {c6288_wire_871, c6288_wire_866});
and_n #(2, 0, 0) AND_522 (c6288_wire_872, {c6288_wire_869_1, c6288_wire_870_1});
and_n #(2, 0, 0) AND_523 (c6288_wire_871, {c6288_wire_873_0, c6288_wire_862_0});
xor_n #(2, 0, 0) XOR_21 (c6288_wire_158, {c6288_wire_874_0, c6288_wire_875_0});
or_n #(2, 0, 0) OR_22 (c6288_wire_874, {c6288_wire_876, c6288_wire_877});
and_n #(2, 0, 0) AND_524 (c6288_wire_878, {c6288_wire_874_1, c6288_wire_875_1});
and_n #(2, 0, 0) AND_525 (c6288_wire_877, {c6288_wire_838, c6288_wire_837_1});
notg #(0, 0) NOT_38 (c6288_wire_876, c6288_wire_879);
xor_n #(2, 0, 0) XOR_22 (c6288_wire_156, {c6288_wire_880_0, c6288_wire_881_0});
or_n #(2, 0, 0) OR_23 (c6288_wire_880, {c6288_wire_878, c6288_wire_882});
and_n #(2, 0, 0) AND_526 (c6288_wire_883, {c6288_wire_880_1, c6288_wire_881_1});
notg #(0, 0) NOT_39 (c6288_wire_882, c6288_wire_884);
xor_n #(2, 0, 0) XOR_23 (c6288_wire_154, {c6288_wire_885_0, c6288_wire_886_0});
or_n #(2, 0, 0) OR_24 (c6288_wire_885, {c6288_wire_883, c6288_wire_887});
and_n #(2, 0, 0) AND_527 (c6288_wire_888, {c6288_wire_885_1, c6288_wire_886_1});
notg #(0, 0) NOT_40 (c6288_wire_887, c6288_wire_889);
xor_n #(2, 0, 0) XOR_24 (c6288_wire_152, {c6288_wire_890_0, c6288_wire_891_0});
or_n #(2, 0, 0) OR_25 (c6288_wire_890, {c6288_wire_888, c6288_wire_892});
and_n #(2, 0, 0) AND_528 (c6288_wire_893, {c6288_wire_890_1, c6288_wire_891_1});
notg #(0, 0) NOT_41 (c6288_wire_892, c6288_wire_894);
xor_n #(2, 0, 0) XOR_25 (c6288_wire_150, {c6288_wire_895_0, c6288_wire_896_0});
or_n #(2, 0, 0) OR_26 (c6288_wire_895, {c6288_wire_893, c6288_wire_897});
and_n #(2, 0, 0) AND_529 (c6288_wire_898, {c6288_wire_895_1, c6288_wire_896_1});
notg #(0, 0) NOT_42 (c6288_wire_897, c6288_wire_899);
xor_n #(2, 0, 0) XOR_26 (c6288_wire_148, {c6288_wire_900_0, c6288_wire_901_0});
or_n #(2, 0, 0) OR_27 (c6288_wire_900, {c6288_wire_898, c6288_wire_902});
and_n #(2, 0, 0) AND_530 (c6288_wire_903, {c6288_wire_900_1, c6288_wire_901_1});
notg #(0, 0) NOT_43 (c6288_wire_902, c6288_wire_904);
xor_n #(2, 0, 0) XOR_27 (c6288_wire_146, {c6288_wire_905_0, c6288_wire_906_0});
or_n #(2, 0, 0) OR_28 (c6288_wire_905, {c6288_wire_903, c6288_wire_907});
and_n #(2, 0, 0) AND_531 (c6288_wire_908, {c6288_wire_905_1, c6288_wire_906_1});
notg #(0, 0) NOT_44 (c6288_wire_907, c6288_wire_909);
xor_n #(2, 0, 0) XOR_28 (c6288_wire_144, {c6288_wire_910_0, c6288_wire_911_0});
or_n #(2, 0, 0) OR_29 (c6288_wire_910, {c6288_wire_908, c6288_wire_912});
and_n #(2, 0, 0) AND_532 (c6288_wire_913, {c6288_wire_910_1, c6288_wire_911_1});
notg #(0, 0) NOT_45 (c6288_wire_912, c6288_wire_914);
xor_n #(2, 0, 0) XOR_29 (c6288_wire_142, {c6288_wire_844_1, c6288_wire_845_1});
or_n #(2, 0, 0) OR_30 (c6288_wire_844, {c6288_wire_913, c6288_wire_915});
notg #(0, 0) NOT_46 (c6288_wire_915, c6288_wire_916);
and_n #(2, 0, 0) AND_533 (c6288_wire_917, {c6288_wire_16_0, c6288_wire_918_0});
notg #(0, 0) NOT_47 (c6288_wire_919, c6288_wire_16_1);
xor_n #(2, 0, 0) XOR_30 (c6288_wire_182, {c6288_wire_920_0, c6288_wire_921_0});
or_n #(2, 0, 0) OR_31 (c6288_wire_920, {c6288_wire_922, c6288_wire_923});
and_n #(2, 0, 0) AND_534 (c6288_wire_924, {c6288_wire_920_1, c6288_wire_921_1});
and_n #(2, 0, 0) AND_535 (c6288_wire_922, {c6288_wire_925_0, c6288_wire_926_0});
notg #(0, 0) NOT_48 (c6288_wire_923, c6288_wire_927);
xor_n #(2, 0, 0) XOR_31 (c6288_wire_180, {c6288_wire_928_0, c6288_wire_929_0});
or_n #(2, 0, 0) OR_32 (c6288_wire_928, {c6288_wire_924, c6288_wire_930});
and_n #(2, 0, 0) AND_536 (c6288_wire_931, {c6288_wire_928_1, c6288_wire_929_1});
notg #(0, 0) NOT_49 (c6288_wire_930, c6288_wire_932);
xor_n #(2, 0, 0) XOR_32 (c6288_wire_178, {c6288_wire_933_0, c6288_wire_934_0});
or_n #(2, 0, 0) OR_33 (c6288_wire_933, {c6288_wire_931, c6288_wire_935});
and_n #(2, 0, 0) AND_537 (c6288_wire_936, {c6288_wire_933_1, c6288_wire_934_1});
notg #(0, 0) NOT_50 (c6288_wire_935, c6288_wire_937);
xor_n #(2, 0, 0) XOR_33 (c6288_wire_176, {c6288_wire_938_0, c6288_wire_939_0});
or_n #(2, 0, 0) OR_34 (c6288_wire_938, {c6288_wire_936, c6288_wire_940});
and_n #(2, 0, 0) AND_538 (c6288_wire_941, {c6288_wire_938_1, c6288_wire_939_1});
notg #(0, 0) NOT_51 (c6288_wire_940, c6288_wire_942);
xor_n #(2, 0, 0) XOR_34 (c6288_wire_870, {c6288_wire_943_0, c6288_wire_944_0});
or_n #(2, 0, 0) OR_35 (c6288_wire_943, {c6288_wire_941, c6288_wire_945});
and_n #(2, 0, 0) AND_539 (c6288_wire_946, {c6288_wire_943_1, c6288_wire_944_1});
notg #(0, 0) NOT_52 (c6288_wire_945, c6288_wire_947);
and_n #(2, 0, 0) AND_540 (c6288_wire_948, {c6288_wire_949_0, c6288_wire_950_0});
or_n #(2, 0, 0) OR_36 (c6288_wire_949, {c6288_wire_872, c6288_wire_946});
and_n #(2, 0, 0) AND_541 (c6288_wire_951, {c6288_wire_949_1, c6288_wire_950_1});
xor_n #(2, 0, 0) XOR_35 (c6288_wire_200, {c6288_wire_952_0, c6288_wire_953_0});
or_n #(2, 0, 0) OR_37 (c6288_wire_952, {c6288_wire_954, c6288_wire_955});
and_n #(2, 0, 0) AND_542 (c6288_wire_956, {c6288_wire_952_1, c6288_wire_953_1});
and_n #(2, 0, 0) AND_543 (c6288_wire_955, {c6288_wire_919, c6288_wire_918_1});
notg #(0, 0) NOT_53 (c6288_wire_954, c6288_wire_957);
xor_n #(2, 0, 0) XOR_36 (c6288_wire_198, {c6288_wire_958_0, c6288_wire_959_0});
or_n #(2, 0, 0) OR_38 (c6288_wire_958, {c6288_wire_956, c6288_wire_960});
and_n #(2, 0, 0) AND_544 (c6288_wire_961, {c6288_wire_958_1, c6288_wire_959_1});
notg #(0, 0) NOT_54 (c6288_wire_960, c6288_wire_962);
xor_n #(2, 0, 0) XOR_37 (c6288_wire_196, {c6288_wire_963_0, c6288_wire_964_0});
or_n #(2, 0, 0) OR_39 (c6288_wire_963, {c6288_wire_961, c6288_wire_965});
and_n #(2, 0, 0) AND_545 (c6288_wire_966, {c6288_wire_963_1, c6288_wire_964_1});
notg #(0, 0) NOT_55 (c6288_wire_965, c6288_wire_967);
xor_n #(2, 0, 0) XOR_38 (c6288_wire_194, {c6288_wire_968_0, c6288_wire_969_0});
or_n #(2, 0, 0) OR_40 (c6288_wire_968, {c6288_wire_966, c6288_wire_970});
and_n #(2, 0, 0) AND_546 (c6288_wire_971, {c6288_wire_968_1, c6288_wire_969_1});
notg #(0, 0) NOT_56 (c6288_wire_970, c6288_wire_972);
xor_n #(2, 0, 0) XOR_39 (c6288_wire_192, {c6288_wire_973_0, c6288_wire_974_0});
or_n #(2, 0, 0) OR_41 (c6288_wire_973, {c6288_wire_971, c6288_wire_975});
and_n #(2, 0, 0) AND_547 (c6288_wire_976, {c6288_wire_973_1, c6288_wire_974_1});
notg #(0, 0) NOT_57 (c6288_wire_975, c6288_wire_977);
xor_n #(2, 0, 0) XOR_40 (c6288_wire_190, {c6288_wire_978_0, c6288_wire_979_0});
or_n #(2, 0, 0) OR_42 (c6288_wire_978, {c6288_wire_976, c6288_wire_980});
and_n #(2, 0, 0) AND_548 (c6288_wire_981, {c6288_wire_978_1, c6288_wire_979_1});
notg #(0, 0) NOT_58 (c6288_wire_980, c6288_wire_982);
xor_n #(2, 0, 0) XOR_41 (c6288_wire_188, {c6288_wire_983_0, c6288_wire_984_0});
or_n #(2, 0, 0) OR_43 (c6288_wire_983, {c6288_wire_981, c6288_wire_985});
and_n #(2, 0, 0) AND_549 (c6288_wire_986, {c6288_wire_983_1, c6288_wire_984_1});
notg #(0, 0) NOT_59 (c6288_wire_985, c6288_wire_987);
xor_n #(2, 0, 0) XOR_42 (c6288_wire_186, {c6288_wire_988_0, c6288_wire_989_0});
or_n #(2, 0, 0) OR_44 (c6288_wire_988, {c6288_wire_986, c6288_wire_990});
and_n #(2, 0, 0) AND_550 (c6288_wire_991, {c6288_wire_988_1, c6288_wire_989_1});
notg #(0, 0) NOT_60 (c6288_wire_990, c6288_wire_992);
xor_n #(2, 0, 0) XOR_43 (c6288_wire_184, {c6288_wire_925_1, c6288_wire_926_1});
or_n #(2, 0, 0) OR_45 (c6288_wire_925, {c6288_wire_991, c6288_wire_993});
notg #(0, 0) NOT_61 (c6288_wire_993, c6288_wire_994);
and_n #(2, 0, 0) AND_551 (c6288_wire_995, {c6288_wire_21_0, c6288_wire_996_0});
notg #(0, 0) NOT_62 (c6288_wire_997, c6288_wire_21_1);
xor_n #(2, 0, 0) XOR_44 (c6288_wire_224, {c6288_wire_998_0, c6288_wire_999_0});
or_n #(2, 0, 0) OR_46 (c6288_wire_998, {c6288_wire_1000, c6288_wire_1001});
and_n #(2, 0, 0) AND_552 (c6288_wire_1002, {c6288_wire_998_1, c6288_wire_999_1});
and_n #(2, 0, 0) AND_553 (c6288_wire_1000, {c6288_wire_1003_0, c6288_wire_1004_0});
notg #(0, 0) NOT_63 (c6288_wire_1001, c6288_wire_1005);
xor_n #(2, 0, 0) XOR_45 (c6288_wire_222, {c6288_wire_1006_0, c6288_wire_1007_0});
or_n #(2, 0, 0) OR_47 (c6288_wire_1006, {c6288_wire_1002, c6288_wire_1008});
and_n #(2, 0, 0) AND_554 (c6288_wire_1009, {c6288_wire_1006_1, c6288_wire_1007_1});
notg #(0, 0) NOT_64 (c6288_wire_1008, c6288_wire_1010);
xor_n #(2, 0, 0) XOR_46 (c6288_wire_220, {c6288_wire_1011_0, c6288_wire_1012_0});
or_n #(2, 0, 0) OR_48 (c6288_wire_1011, {c6288_wire_1009, c6288_wire_1013});
and_n #(2, 0, 0) AND_555 (c6288_wire_1014, {c6288_wire_1011_1, c6288_wire_1012_1});
notg #(0, 0) NOT_65 (c6288_wire_1013, c6288_wire_1015);
xor_n #(2, 0, 0) XOR_47 (c6288_wire_218, {c6288_wire_1016_0, c6288_wire_1017_0});
or_n #(2, 0, 0) OR_49 (c6288_wire_1016, {c6288_wire_1014, c6288_wire_1018});
and_n #(2, 0, 0) AND_556 (c6288_wire_1019, {c6288_wire_1016_1, c6288_wire_1017_1});
notg #(0, 0) NOT_66 (c6288_wire_1018, c6288_wire_1020);
xor_n #(2, 0, 0) XOR_48 (c6288_wire_950, {c6288_wire_1021_0, c6288_wire_1022_0});
or_n #(2, 0, 0) OR_50 (c6288_wire_1021, {c6288_wire_1019, c6288_wire_1023});
and_n #(2, 0, 0) AND_557 (c6288_wire_1024, {c6288_wire_1021_1, c6288_wire_1022_1});
notg #(0, 0) NOT_67 (c6288_wire_1023, c6288_wire_1025);
and_n #(2, 0, 0) AND_558 (c6288_wire_1026, {c6288_wire_1027_0, c6288_wire_1028_0});
or_n #(2, 0, 0) OR_51 (c6288_wire_1027, {c6288_wire_951, c6288_wire_1024});
and_n #(2, 0, 0) AND_559 (c6288_wire_1029, {c6288_wire_1027_1, c6288_wire_1028_1});
xor_n #(2, 0, 0) XOR_49 (c6288_wire_242, {c6288_wire_1030_0, c6288_wire_1031_0});
or_n #(2, 0, 0) OR_52 (c6288_wire_1030, {c6288_wire_1032, c6288_wire_1033});
and_n #(2, 0, 0) AND_560 (c6288_wire_1034, {c6288_wire_1030_1, c6288_wire_1031_1});
and_n #(2, 0, 0) AND_561 (c6288_wire_1033, {c6288_wire_997, c6288_wire_996_1});
notg #(0, 0) NOT_68 (c6288_wire_1032, c6288_wire_1035);
xor_n #(2, 0, 0) XOR_50 (c6288_wire_240, {c6288_wire_1036_0, c6288_wire_1037_0});
or_n #(2, 0, 0) OR_53 (c6288_wire_1036, {c6288_wire_1034, c6288_wire_1038});
and_n #(2, 0, 0) AND_562 (c6288_wire_1039, {c6288_wire_1036_1, c6288_wire_1037_1});
notg #(0, 0) NOT_69 (c6288_wire_1038, c6288_wire_1040);
xor_n #(2, 0, 0) XOR_51 (c6288_wire_238, {c6288_wire_1041_0, c6288_wire_1042_0});
or_n #(2, 0, 0) OR_54 (c6288_wire_1041, {c6288_wire_1039, c6288_wire_1043});
and_n #(2, 0, 0) AND_563 (c6288_wire_1044, {c6288_wire_1041_1, c6288_wire_1042_1});
notg #(0, 0) NOT_70 (c6288_wire_1043, c6288_wire_1045);
xor_n #(2, 0, 0) XOR_52 (c6288_wire_236, {c6288_wire_1046_0, c6288_wire_1047_0});
or_n #(2, 0, 0) OR_55 (c6288_wire_1046, {c6288_wire_1044, c6288_wire_1048});
and_n #(2, 0, 0) AND_564 (c6288_wire_1049, {c6288_wire_1046_1, c6288_wire_1047_1});
notg #(0, 0) NOT_71 (c6288_wire_1048, c6288_wire_1050);
xor_n #(2, 0, 0) XOR_53 (c6288_wire_234, {c6288_wire_1051_0, c6288_wire_1052_0});
or_n #(2, 0, 0) OR_56 (c6288_wire_1051, {c6288_wire_1049, c6288_wire_1053});
and_n #(2, 0, 0) AND_565 (c6288_wire_1054, {c6288_wire_1051_1, c6288_wire_1052_1});
notg #(0, 0) NOT_72 (c6288_wire_1053, c6288_wire_1055);
xor_n #(2, 0, 0) XOR_54 (c6288_wire_232, {c6288_wire_1056_0, c6288_wire_1057_0});
or_n #(2, 0, 0) OR_57 (c6288_wire_1056, {c6288_wire_1054, c6288_wire_1058});
and_n #(2, 0, 0) AND_566 (c6288_wire_1059, {c6288_wire_1056_1, c6288_wire_1057_1});
notg #(0, 0) NOT_73 (c6288_wire_1058, c6288_wire_1060);
xor_n #(2, 0, 0) XOR_55 (c6288_wire_230, {c6288_wire_1061_0, c6288_wire_1062_0});
or_n #(2, 0, 0) OR_58 (c6288_wire_1061, {c6288_wire_1059, c6288_wire_1063});
and_n #(2, 0, 0) AND_567 (c6288_wire_1064, {c6288_wire_1061_1, c6288_wire_1062_1});
notg #(0, 0) NOT_74 (c6288_wire_1063, c6288_wire_1065);
xor_n #(2, 0, 0) XOR_56 (c6288_wire_228, {c6288_wire_1066_0, c6288_wire_1067_0});
or_n #(2, 0, 0) OR_59 (c6288_wire_1066, {c6288_wire_1064, c6288_wire_1068});
and_n #(2, 0, 0) AND_568 (c6288_wire_1069, {c6288_wire_1066_1, c6288_wire_1067_1});
notg #(0, 0) NOT_75 (c6288_wire_1068, c6288_wire_1070);
xor_n #(2, 0, 0) XOR_57 (c6288_wire_226, {c6288_wire_1003_1, c6288_wire_1004_1});
or_n #(2, 0, 0) OR_60 (c6288_wire_1003, {c6288_wire_1069, c6288_wire_1071});
notg #(0, 0) NOT_76 (c6288_wire_1071, c6288_wire_1072);
xor_n #(2, 0, 0) XOR_58 (c6288_wire_286, {c6288_wire_26_0, c6288_wire_1073_0});
xor_n #(2, 0, 0) XOR_59 (c6288_wire_266, {c6288_wire_1074_0, c6288_wire_1075_0});
or_n #(2, 0, 0) OR_61 (c6288_wire_1074, {c6288_wire_1076, c6288_wire_1077});
and_n #(2, 0, 0) AND_569 (c6288_wire_1078, {c6288_wire_1074_1, c6288_wire_1075_1});
and_n #(2, 0, 0) AND_570 (c6288_wire_1076, {c6288_wire_1079_0, c6288_wire_1080_0});
notg #(0, 0) NOT_77 (c6288_wire_1077, c6288_wire_1081);
xor_n #(2, 0, 0) XOR_60 (c6288_wire_264, {c6288_wire_1082_0, c6288_wire_1083_0});
or_n #(2, 0, 0) OR_62 (c6288_wire_1082, {c6288_wire_1078, c6288_wire_1084});
and_n #(2, 0, 0) AND_571 (c6288_wire_1085, {c6288_wire_1082_1, c6288_wire_1083_1});
notg #(0, 0) NOT_78 (c6288_wire_1084, c6288_wire_1086);
xor_n #(2, 0, 0) XOR_61 (c6288_wire_262, {c6288_wire_1087_0, c6288_wire_1088_0});
or_n #(2, 0, 0) OR_63 (c6288_wire_1087, {c6288_wire_1085, c6288_wire_1089});
and_n #(2, 0, 0) AND_572 (c6288_wire_1090, {c6288_wire_1087_1, c6288_wire_1088_1});
notg #(0, 0) NOT_79 (c6288_wire_1089, c6288_wire_1091);
xor_n #(2, 0, 0) XOR_62 (c6288_wire_260, {c6288_wire_1092_0, c6288_wire_1093_0});
or_n #(2, 0, 0) OR_64 (c6288_wire_1092, {c6288_wire_1090, c6288_wire_1094});
and_n #(2, 0, 0) AND_573 (c6288_wire_1095, {c6288_wire_1092_1, c6288_wire_1093_1});
notg #(0, 0) NOT_80 (c6288_wire_1094, c6288_wire_1096);
xor_n #(2, 0, 0) XOR_63 (c6288_wire_1028, {c6288_wire_1097_0, c6288_wire_1098_0});
or_n #(2, 0, 0) OR_65 (c6288_wire_1097, {c6288_wire_1095, c6288_wire_1099});
and_n #(2, 0, 0) AND_574 (c6288_wire_1100, {c6288_wire_1097_1, c6288_wire_1098_1});
notg #(0, 0) NOT_81 (c6288_wire_1099, c6288_wire_1101);
and_n #(2, 0, 0) AND_575 (c6288_wire_1102, {c6288_wire_1103_0, c6288_wire_1104_0});
or_n #(2, 0, 0) OR_66 (c6288_wire_1103, {c6288_wire_1029, c6288_wire_1100});
notg #(0, 0) NOT_82 (c6288_wire_1105, c6288_wire_1103_1);
notg #(0, 0) NOT_83 (c6288_wire_1106, c6288_wire_1103_2);
and_n #(2, 0, 0) AND_576 (c6288_wire_1107, {c6288_wire_1108_0, c6288_wire_1109_0});
or_n #(2, 0, 0) OR_67 (c6288_wire_1108, {c6288_wire_1110, c6288_wire_1111});
and_n #(2, 0, 0) AND_577 (c6288_wire_1112, {c6288_wire_1108_1, c6288_wire_1113});
nor_n #(2, 0, 0) NOR_2 (c6288_wire_1111, {c6288_wire_26_1, c6288_wire_1073_1});
notg #(0, 0) NOT_84 (c6288_wire_1110, c6288_wire_1114);
xor_n #(2, 0, 0) XOR_64 (c6288_wire_282, {c6288_wire_1115_0, c6288_wire_1116_0});
or_n #(2, 0, 0) OR_68 (c6288_wire_1115, {c6288_wire_1117, c6288_wire_1112});
and_n #(2, 0, 0) AND_578 (c6288_wire_1118, {c6288_wire_1115_1, c6288_wire_1116_1});
notg #(0, 0) NOT_85 (c6288_wire_1113, c6288_wire_1109_1);
notg #(0, 0) NOT_86 (c6288_wire_1117, c6288_wire_1119);
xor_n #(2, 0, 0) XOR_65 (c6288_wire_280, {c6288_wire_1120_0, c6288_wire_1121_0});
or_n #(2, 0, 0) OR_69 (c6288_wire_1120, {c6288_wire_1118, c6288_wire_1122});
and_n #(2, 0, 0) AND_579 (c6288_wire_1123, {c6288_wire_1120_1, c6288_wire_1121_1});
notg #(0, 0) NOT_87 (c6288_wire_1122, c6288_wire_1124);
xor_n #(2, 0, 0) XOR_66 (c6288_wire_278, {c6288_wire_1125_0, c6288_wire_1126_0});
or_n #(2, 0, 0) OR_70 (c6288_wire_1125, {c6288_wire_1123, c6288_wire_1127});
and_n #(2, 0, 0) AND_580 (c6288_wire_1128, {c6288_wire_1125_1, c6288_wire_1126_1});
notg #(0, 0) NOT_88 (c6288_wire_1127, c6288_wire_1129);
xor_n #(2, 0, 0) XOR_67 (c6288_wire_276, {c6288_wire_1130_0, c6288_wire_1131_0});
or_n #(2, 0, 0) OR_71 (c6288_wire_1130, {c6288_wire_1128, c6288_wire_1132});
and_n #(2, 0, 0) AND_581 (c6288_wire_1133, {c6288_wire_1130_1, c6288_wire_1131_1});
notg #(0, 0) NOT_89 (c6288_wire_1132, c6288_wire_1134);
xor_n #(2, 0, 0) XOR_68 (c6288_wire_274, {c6288_wire_1135_0, c6288_wire_1136_0});
or_n #(2, 0, 0) OR_72 (c6288_wire_1135, {c6288_wire_1133, c6288_wire_1137});
and_n #(2, 0, 0) AND_582 (c6288_wire_1138, {c6288_wire_1135_1, c6288_wire_1136_1});
notg #(0, 0) NOT_90 (c6288_wire_1137, c6288_wire_1139);
xor_n #(2, 0, 0) XOR_69 (c6288_wire_272, {c6288_wire_1140_0, c6288_wire_1141_0});
or_n #(2, 0, 0) OR_73 (c6288_wire_1140, {c6288_wire_1138, c6288_wire_1142});
and_n #(2, 0, 0) AND_583 (c6288_wire_1143, {c6288_wire_1140_1, c6288_wire_1141_1});
notg #(0, 0) NOT_91 (c6288_wire_1142, c6288_wire_1144);
xor_n #(2, 0, 0) XOR_70 (c6288_wire_270, {c6288_wire_1145_0, c6288_wire_1146_0});
or_n #(2, 0, 0) OR_74 (c6288_wire_1145, {c6288_wire_1143, c6288_wire_1147});
and_n #(2, 0, 0) AND_584 (c6288_wire_1148, {c6288_wire_1145_1, c6288_wire_1146_1});
notg #(0, 0) NOT_92 (c6288_wire_1147, c6288_wire_1149);
xor_n #(2, 0, 0) XOR_71 (c6288_wire_268, {c6288_wire_1079_1, c6288_wire_1080_1});
or_n #(2, 0, 0) OR_75 (c6288_wire_1079, {c6288_wire_1148, c6288_wire_1150});
notg #(0, 0) NOT_93 (c6288_wire_1150, c6288_wire_1151);
and_n #(2, 0, 0) AND_585 (c6288_wire_1152, {c6288_wire_1153, c6288_wire_1154});
or_n #(2, 0, 0) OR_76 (c6288_wire_1155, {c6288_wire_1152_0, c6288_wire_338});
notg #(0, 0) NOT_94 (c6288_wire_1156, c6288_wire_1152_1);
and_n #(2, 0, 0) AND_586 (c6288_wire_1157, {c6288_wire_1152_2, c6288_wire_1158});
and_n #(2, 0, 0) AND_587 (c6288_wire_1159, {c6288_wire_1155, c6288_wire_1160});
or_n #(2, 0, 0) OR_77 (c6288_wire_1161, {c6288_wire_1159_0, c6288_wire_339});
notg #(0, 0) NOT_95 (c6288_wire_1162, c6288_wire_1159_1);
and_n #(2, 0, 0) AND_588 (c6288_wire_1163, {c6288_wire_1159_2, c6288_wire_1164});
and_n #(2, 0, 0) AND_589 (c6288_wire_1165, {c6288_wire_1161, c6288_wire_1166});
or_n #(2, 0, 0) OR_78 (c6288_wire_1167, {c6288_wire_1165_0, c6288_wire_340});
notg #(0, 0) NOT_96 (c6288_wire_1168, c6288_wire_1165_1);
and_n #(2, 0, 0) AND_590 (c6288_wire_1169, {c6288_wire_1165_2, c6288_wire_1170});
and_n #(2, 0, 0) AND_591 (c6288_wire_1171, {c6288_wire_1167, c6288_wire_1172});
or_n #(2, 0, 0) OR_79 (c6288_wire_1173, {c6288_wire_1171_0, c6288_wire_341});
notg #(0, 0) NOT_97 (c6288_wire_1174, c6288_wire_1171_1);
and_n #(2, 0, 0) AND_592 (c6288_wire_1175, {c6288_wire_1171_2, c6288_wire_1176});
and_n #(2, 0, 0) AND_593 (c6288_wire_1177, {c6288_wire_1173, c6288_wire_1178});
notg #(0, 0) NOT_98 (c6288_wire_1179, c6288_wire_1177_0);
and_n #(2, 0, 0) AND_594 (c6288_wire_1180, {c6288_wire_1177_1, c6288_wire_1181});
and_n #(2, 0, 0) AND_595 (c6288_wire_1182, {c6288_wire_1177_2, c6288_wire_1105});
or_n #(2, 0, 0) OR_80 (c6288_wire_1183, {c6288_wire_1177_3, c6288_wire_1106});
and_n #(2, 0, 0) AND_596 (c6288_wire_1184, {c6288_wire_357, c6288_wire_1183});
or_n #(2, 0, 0) OR_81 (c6288_wire_1185, {c6288_wire_1182, c6288_wire_1184});
and_n #(2, 0, 0) AND_597 (c6288_wire_1186, {c6288_wire_358, c6288_wire_1187});
or_n #(2, 0, 0) OR_82 (c6288_wire_1188, {c6288_wire_1186_0, c6288_wire_329});
notg #(0, 0) NOT_99 (c6288_wire_1189, c6288_wire_1186_1);
and_n #(2, 0, 0) AND_598 (c6288_wire_1190, {c6288_wire_1186_2, c6288_wire_1191});
and_n #(2, 0, 0) AND_599 (c6288_wire_1192, {c6288_wire_1188, c6288_wire_1193});
or_n #(2, 0, 0) OR_83 (c6288_wire_1194, {c6288_wire_1192_0, c6288_wire_331});
notg #(0, 0) NOT_100 (c6288_wire_1195, c6288_wire_1192_1);
and_n #(2, 0, 0) AND_600 (c6288_wire_1196, {c6288_wire_1192_2, c6288_wire_1197});
and_n #(2, 0, 0) AND_601 (c6288_wire_1198, {c6288_wire_1194, c6288_wire_1199});
or_n #(2, 0, 0) OR_84 (c6288_wire_1200, {c6288_wire_1198_0, c6288_wire_332});
notg #(0, 0) NOT_101 (c6288_wire_1201, c6288_wire_1198_1);
and_n #(2, 0, 0) AND_602 (c6288_wire_1202, {c6288_wire_1198_2, c6288_wire_1203});
and_n #(2, 0, 0) AND_603 (c6288_wire_1204, {c6288_wire_1200, c6288_wire_1205});
or_n #(2, 0, 0) OR_85 (c6288_wire_1206, {c6288_wire_1204_0, c6288_wire_333});
notg #(0, 0) NOT_102 (c6288_wire_1207, c6288_wire_1204_1);
and_n #(2, 0, 0) AND_604 (c6288_wire_1208, {c6288_wire_1204_2, c6288_wire_1209});
and_n #(2, 0, 0) AND_605 (c6288_wire_1210, {c6288_wire_1206, c6288_wire_1211});
or_n #(2, 0, 0) OR_86 (c6288_wire_1212, {c6288_wire_1210_0, c6288_wire_334});
notg #(0, 0) NOT_103 (c6288_wire_1213, c6288_wire_1210_1);
and_n #(2, 0, 0) AND_606 (c6288_wire_1214, {c6288_wire_1210_2, c6288_wire_1215});
and_n #(2, 0, 0) AND_607 (c6288_wire_1216, {c6288_wire_1212, c6288_wire_1217});
or_n #(2, 0, 0) OR_87 (c6288_wire_1218, {c6288_wire_1216_0, c6288_wire_335});
notg #(0, 0) NOT_104 (c6288_wire_1219, c6288_wire_1216_1);
and_n #(2, 0, 0) AND_608 (c6288_wire_1220, {c6288_wire_1216_2, c6288_wire_1221});
and_n #(2, 0, 0) AND_609 (c6288_wire_1222, {c6288_wire_1218, c6288_wire_1223});
or_n #(2, 0, 0) OR_88 (c6288_wire_1224, {c6288_wire_1222_0, c6288_wire_336});
notg #(0, 0) NOT_105 (c6288_wire_1225, c6288_wire_1222_1);
and_n #(2, 0, 0) AND_610 (c6288_wire_1226, {c6288_wire_1222_2, c6288_wire_1227});
and_n #(2, 0, 0) AND_611 (c6288_wire_1228, {c6288_wire_1224, c6288_wire_1229});
or_n #(2, 0, 0) OR_89 (c6288_wire_1153, {c6288_wire_1228_0, c6288_wire_337});
notg #(0, 0) NOT_106 (c6288_wire_1230, c6288_wire_1228_1);
and_n #(2, 0, 0) AND_612 (c6288_wire_1231, {c6288_wire_1228_2, c6288_wire_1232});
and_n #(2, 0, 0) AND_613 (c6288_wire_1233, {c6288_wire_38_0, c6288_wire_1234_0});
notg #(0, 0) NOT_107 (c6288_wire_1235, c6288_wire_38_1);
xor_n #(2, 0, 0) XOR_72 (c6288_wire_382, {c6288_wire_1236_0, c6288_wire_1237_0});
or_n #(2, 0, 0) OR_90 (c6288_wire_1236, {c6288_wire_1238, c6288_wire_1239});
and_n #(2, 0, 0) AND_614 (c6288_wire_1240, {c6288_wire_1236_1, c6288_wire_1237_1});
and_n #(2, 0, 0) AND_615 (c6288_wire_1238, {c6288_wire_1241_0, c6288_wire_1242_0});
notg #(0, 0) NOT_108 (c6288_wire_1239, c6288_wire_1243);
xor_n #(2, 0, 0) XOR_73 (c6288_wire_380, {c6288_wire_1244_0, c6288_wire_1245_0});
or_n #(2, 0, 0) OR_91 (c6288_wire_1244, {c6288_wire_1240, c6288_wire_1246});
and_n #(2, 0, 0) AND_616 (c6288_wire_1247, {c6288_wire_1244_1, c6288_wire_1245_1});
notg #(0, 0) NOT_109 (c6288_wire_1246, c6288_wire_1248);
xor_n #(2, 0, 0) XOR_74 (c6288_wire_378, {c6288_wire_1249_0, c6288_wire_1250_0});
or_n #(2, 0, 0) OR_92 (c6288_wire_1249, {c6288_wire_1247, c6288_wire_1251});
and_n #(2, 0, 0) AND_617 (c6288_wire_1252, {c6288_wire_1249_1, c6288_wire_1250_1});
notg #(0, 0) NOT_110 (c6288_wire_1251, c6288_wire_1253);
xor_n #(2, 0, 0) XOR_75 (c6288_wire_376, {c6288_wire_1254_0, c6288_wire_1255_0});
or_n #(2, 0, 0) OR_93 (c6288_wire_1254, {c6288_wire_1252, c6288_wire_1256});
and_n #(2, 0, 0) AND_618 (c6288_wire_1257, {c6288_wire_1254_1, c6288_wire_1255_1});
notg #(0, 0) NOT_111 (c6288_wire_1256, c6288_wire_1258);
xor_n #(2, 0, 0) XOR_76 (c6288_wire_782, {c6288_wire_1259_0, c6288_wire_1260_0});
or_n #(2, 0, 0) OR_94 (c6288_wire_1259, {c6288_wire_1257, c6288_wire_1261});
and_n #(2, 0, 0) AND_619 (c6288_wire_1262, {c6288_wire_1259_1, c6288_wire_1260_1});
notg #(0, 0) NOT_112 (c6288_wire_1261, c6288_wire_1263);
and_n #(2, 0, 0) AND_620 (c6288_wire_1264, {c6288_wire_1265_0, c6288_wire_1266_0});
and_n #(2, 0, 0) AND_621 (c6288_wire_1267, {c6288_wire_1265_1, c6288_wire_1266_1});
or_n #(2, 0, 0) OR_95 (c6288_wire_1265, {c6288_wire_1262, c6288_wire_1268});
and_n #(2, 0, 0) AND_622 (c6288_wire_1268, {c6288_wire_783, c6288_wire_782_1});
xor_n #(2, 0, 0) XOR_77 (c6288_wire_400, {c6288_wire_1269_0, c6288_wire_1270_0});
or_n #(2, 0, 0) OR_96 (c6288_wire_1269, {c6288_wire_1271, c6288_wire_1272});
and_n #(2, 0, 0) AND_623 (c6288_wire_1273, {c6288_wire_1269_1, c6288_wire_1270_1});
and_n #(2, 0, 0) AND_624 (c6288_wire_1272, {c6288_wire_1235, c6288_wire_1234_1});
notg #(0, 0) NOT_113 (c6288_wire_1271, c6288_wire_1274);
xor_n #(2, 0, 0) XOR_78 (c6288_wire_398, {c6288_wire_1275_0, c6288_wire_1276_0});
or_n #(2, 0, 0) OR_97 (c6288_wire_1275, {c6288_wire_1273, c6288_wire_1277});
and_n #(2, 0, 0) AND_625 (c6288_wire_1278, {c6288_wire_1275_1, c6288_wire_1276_1});
notg #(0, 0) NOT_114 (c6288_wire_1277, c6288_wire_1279);
xor_n #(2, 0, 0) XOR_79 (c6288_wire_396, {c6288_wire_1280_0, c6288_wire_1281_0});
or_n #(2, 0, 0) OR_98 (c6288_wire_1280, {c6288_wire_1278, c6288_wire_1282});
and_n #(2, 0, 0) AND_626 (c6288_wire_1283, {c6288_wire_1280_1, c6288_wire_1281_1});
notg #(0, 0) NOT_115 (c6288_wire_1282, c6288_wire_1284);
xor_n #(2, 0, 0) XOR_80 (c6288_wire_394, {c6288_wire_1285_0, c6288_wire_1286_0});
or_n #(2, 0, 0) OR_99 (c6288_wire_1285, {c6288_wire_1283, c6288_wire_1287});
and_n #(2, 0, 0) AND_627 (c6288_wire_1288, {c6288_wire_1285_1, c6288_wire_1286_1});
notg #(0, 0) NOT_116 (c6288_wire_1287, c6288_wire_1289);
xor_n #(2, 0, 0) XOR_81 (c6288_wire_392, {c6288_wire_1290_0, c6288_wire_1291_0});
or_n #(2, 0, 0) OR_100 (c6288_wire_1290, {c6288_wire_1288, c6288_wire_1292});
and_n #(2, 0, 0) AND_628 (c6288_wire_1293, {c6288_wire_1290_1, c6288_wire_1291_1});
notg #(0, 0) NOT_117 (c6288_wire_1292, c6288_wire_1294);
xor_n #(2, 0, 0) XOR_82 (c6288_wire_390, {c6288_wire_1295_0, c6288_wire_1296_0});
or_n #(2, 0, 0) OR_101 (c6288_wire_1295, {c6288_wire_1293, c6288_wire_1297});
and_n #(2, 0, 0) AND_629 (c6288_wire_1298, {c6288_wire_1295_1, c6288_wire_1296_1});
notg #(0, 0) NOT_118 (c6288_wire_1297, c6288_wire_1299);
xor_n #(2, 0, 0) XOR_83 (c6288_wire_388, {c6288_wire_1300_0, c6288_wire_1301_0});
or_n #(2, 0, 0) OR_102 (c6288_wire_1300, {c6288_wire_1298, c6288_wire_1302});
and_n #(2, 0, 0) AND_630 (c6288_wire_1303, {c6288_wire_1300_1, c6288_wire_1301_1});
notg #(0, 0) NOT_119 (c6288_wire_1302, c6288_wire_1304);
xor_n #(2, 0, 0) XOR_84 (c6288_wire_386, {c6288_wire_1305_0, c6288_wire_1306_0});
or_n #(2, 0, 0) OR_103 (c6288_wire_1305, {c6288_wire_1303, c6288_wire_1307});
and_n #(2, 0, 0) AND_631 (c6288_wire_1308, {c6288_wire_1305_1, c6288_wire_1306_1});
notg #(0, 0) NOT_120 (c6288_wire_1307, c6288_wire_1309);
xor_n #(2, 0, 0) XOR_85 (c6288_wire_384, {c6288_wire_1241_1, c6288_wire_1242_1});
or_n #(2, 0, 0) OR_104 (c6288_wire_1241, {c6288_wire_1308, c6288_wire_1310});
notg #(0, 0) NOT_121 (c6288_wire_1310, c6288_wire_1311);
and_n #(2, 0, 0) AND_632 (c6288_wire_1312, {c6288_wire_43_0, c6288_wire_1313_0});
notg #(0, 0) NOT_122 (c6288_wire_1314, c6288_wire_43_1);
xor_n #(2, 0, 0) XOR_86 (c6288_wire_424, {c6288_wire_1315_0, c6288_wire_1316_0});
or_n #(2, 0, 0) OR_105 (c6288_wire_1315, {c6288_wire_1317, c6288_wire_1318});
and_n #(2, 0, 0) AND_633 (c6288_wire_1319, {c6288_wire_1315_1, c6288_wire_1316_1});
and_n #(2, 0, 0) AND_634 (c6288_wire_1317, {c6288_wire_1320_0, c6288_wire_1321_0});
notg #(0, 0) NOT_123 (c6288_wire_1318, c6288_wire_1322);
xor_n #(2, 0, 0) XOR_87 (c6288_wire_422, {c6288_wire_1323_0, c6288_wire_1324_0});
or_n #(2, 0, 0) OR_106 (c6288_wire_1323, {c6288_wire_1319, c6288_wire_1325});
and_n #(2, 0, 0) AND_635 (c6288_wire_1326, {c6288_wire_1323_1, c6288_wire_1324_1});
notg #(0, 0) NOT_124 (c6288_wire_1325, c6288_wire_1327);
xor_n #(2, 0, 0) XOR_88 (c6288_wire_420, {c6288_wire_1328_0, c6288_wire_1329_0});
or_n #(2, 0, 0) OR_107 (c6288_wire_1328, {c6288_wire_1326, c6288_wire_1330});
and_n #(2, 0, 0) AND_636 (c6288_wire_1331, {c6288_wire_1328_1, c6288_wire_1329_1});
notg #(0, 0) NOT_125 (c6288_wire_1330, c6288_wire_1332);
xor_n #(2, 0, 0) XOR_89 (c6288_wire_418, {c6288_wire_1333_0, c6288_wire_1334_0});
or_n #(2, 0, 0) OR_108 (c6288_wire_1333, {c6288_wire_1331, c6288_wire_1335});
and_n #(2, 0, 0) AND_637 (c6288_wire_1336, {c6288_wire_1333_1, c6288_wire_1334_1});
notg #(0, 0) NOT_126 (c6288_wire_1335, c6288_wire_1337);
xor_n #(2, 0, 0) XOR_90 (c6288_wire_1266, {c6288_wire_1338_0, c6288_wire_1339_0});
or_n #(2, 0, 0) OR_109 (c6288_wire_1338, {c6288_wire_1336, c6288_wire_1340});
and_n #(2, 0, 0) AND_638 (c6288_wire_1341, {c6288_wire_1338_1, c6288_wire_1339_1});
notg #(0, 0) NOT_127 (c6288_wire_1340, c6288_wire_1342);
and_n #(2, 0, 0) AND_639 (c6288_wire_1343, {c6288_wire_1344_0, c6288_wire_1345_0});
or_n #(2, 0, 0) OR_110 (c6288_wire_1344, {c6288_wire_1267, c6288_wire_1341});
and_n #(2, 0, 0) AND_640 (c6288_wire_1346, {c6288_wire_1344_1, c6288_wire_1345_1});
xor_n #(2, 0, 0) XOR_91 (c6288_wire_442, {c6288_wire_1347_0, c6288_wire_1348_0});
or_n #(2, 0, 0) OR_111 (c6288_wire_1347, {c6288_wire_1349, c6288_wire_1350});
and_n #(2, 0, 0) AND_641 (c6288_wire_1351, {c6288_wire_1347_1, c6288_wire_1348_1});
and_n #(2, 0, 0) AND_642 (c6288_wire_1350, {c6288_wire_1314, c6288_wire_1313_1});
notg #(0, 0) NOT_128 (c6288_wire_1349, c6288_wire_1352);
xor_n #(2, 0, 0) XOR_92 (c6288_wire_440, {c6288_wire_1353_0, c6288_wire_1354_0});
or_n #(2, 0, 0) OR_112 (c6288_wire_1353, {c6288_wire_1351, c6288_wire_1355});
and_n #(2, 0, 0) AND_643 (c6288_wire_1356, {c6288_wire_1353_1, c6288_wire_1354_1});
notg #(0, 0) NOT_129 (c6288_wire_1355, c6288_wire_1357);
xor_n #(2, 0, 0) XOR_93 (c6288_wire_438, {c6288_wire_1358_0, c6288_wire_1359_0});
or_n #(2, 0, 0) OR_113 (c6288_wire_1358, {c6288_wire_1356, c6288_wire_1360});
and_n #(2, 0, 0) AND_644 (c6288_wire_1361, {c6288_wire_1358_1, c6288_wire_1359_1});
notg #(0, 0) NOT_130 (c6288_wire_1360, c6288_wire_1362);
xor_n #(2, 0, 0) XOR_94 (c6288_wire_436, {c6288_wire_1363_0, c6288_wire_1364_0});
or_n #(2, 0, 0) OR_114 (c6288_wire_1363, {c6288_wire_1361, c6288_wire_1365});
and_n #(2, 0, 0) AND_645 (c6288_wire_1366, {c6288_wire_1363_1, c6288_wire_1364_1});
notg #(0, 0) NOT_131 (c6288_wire_1365, c6288_wire_1367);
xor_n #(2, 0, 0) XOR_95 (c6288_wire_434, {c6288_wire_1368_0, c6288_wire_1369_0});
or_n #(2, 0, 0) OR_115 (c6288_wire_1368, {c6288_wire_1366, c6288_wire_1370});
and_n #(2, 0, 0) AND_646 (c6288_wire_1371, {c6288_wire_1368_1, c6288_wire_1369_1});
notg #(0, 0) NOT_132 (c6288_wire_1370, c6288_wire_1372);
xor_n #(2, 0, 0) XOR_96 (c6288_wire_432, {c6288_wire_1373_0, c6288_wire_1374_0});
or_n #(2, 0, 0) OR_116 (c6288_wire_1373, {c6288_wire_1371, c6288_wire_1375});
and_n #(2, 0, 0) AND_647 (c6288_wire_1376, {c6288_wire_1373_1, c6288_wire_1374_1});
notg #(0, 0) NOT_133 (c6288_wire_1375, c6288_wire_1377);
xor_n #(2, 0, 0) XOR_97 (c6288_wire_430, {c6288_wire_1378_0, c6288_wire_1379_0});
or_n #(2, 0, 0) OR_117 (c6288_wire_1378, {c6288_wire_1376, c6288_wire_1380});
and_n #(2, 0, 0) AND_648 (c6288_wire_1381, {c6288_wire_1378_1, c6288_wire_1379_1});
notg #(0, 0) NOT_134 (c6288_wire_1380, c6288_wire_1382);
xor_n #(2, 0, 0) XOR_98 (c6288_wire_428, {c6288_wire_1383_0, c6288_wire_1384_0});
or_n #(2, 0, 0) OR_118 (c6288_wire_1383, {c6288_wire_1381, c6288_wire_1385});
and_n #(2, 0, 0) AND_649 (c6288_wire_1386, {c6288_wire_1383_1, c6288_wire_1384_1});
notg #(0, 0) NOT_135 (c6288_wire_1385, c6288_wire_1387);
xor_n #(2, 0, 0) XOR_99 (c6288_wire_426, {c6288_wire_1320_1, c6288_wire_1321_1});
or_n #(2, 0, 0) OR_119 (c6288_wire_1320, {c6288_wire_1386, c6288_wire_1388});
notg #(0, 0) NOT_136 (c6288_wire_1388, c6288_wire_1389);
and_n #(2, 0, 0) AND_650 (c6288_wire_1390, {c6288_wire_48_0, c6288_wire_1391_0});
notg #(0, 0) NOT_137 (c6288_wire_1392, c6288_wire_48_1);
xor_n #(2, 0, 0) XOR_100 (c6288_wire_466, {c6288_wire_1393_0, c6288_wire_1394_0});
or_n #(2, 0, 0) OR_120 (c6288_wire_1393, {c6288_wire_1395, c6288_wire_1396});
and_n #(2, 0, 0) AND_651 (c6288_wire_1397, {c6288_wire_1393_1, c6288_wire_1394_1});
and_n #(2, 0, 0) AND_652 (c6288_wire_1395, {c6288_wire_1398_0, c6288_wire_1399_0});
notg #(0, 0) NOT_138 (c6288_wire_1396, c6288_wire_1400);
xor_n #(2, 0, 0) XOR_101 (c6288_wire_464, {c6288_wire_1401_0, c6288_wire_1402_0});
or_n #(2, 0, 0) OR_121 (c6288_wire_1401, {c6288_wire_1397, c6288_wire_1403});
and_n #(2, 0, 0) AND_653 (c6288_wire_1404, {c6288_wire_1401_1, c6288_wire_1402_1});
notg #(0, 0) NOT_139 (c6288_wire_1403, c6288_wire_1405);
xor_n #(2, 0, 0) XOR_102 (c6288_wire_462, {c6288_wire_1406_0, c6288_wire_1407_0});
or_n #(2, 0, 0) OR_122 (c6288_wire_1406, {c6288_wire_1404, c6288_wire_1408});
and_n #(2, 0, 0) AND_654 (c6288_wire_1409, {c6288_wire_1406_1, c6288_wire_1407_1});
notg #(0, 0) NOT_140 (c6288_wire_1408, c6288_wire_1410);
xor_n #(2, 0, 0) XOR_103 (c6288_wire_460, {c6288_wire_1411_0, c6288_wire_1412_0});
or_n #(2, 0, 0) OR_123 (c6288_wire_1411, {c6288_wire_1409, c6288_wire_1413});
and_n #(2, 0, 0) AND_655 (c6288_wire_1414, {c6288_wire_1411_1, c6288_wire_1412_1});
notg #(0, 0) NOT_141 (c6288_wire_1413, c6288_wire_1415);
xor_n #(2, 0, 0) XOR_104 (c6288_wire_1345, {c6288_wire_1416_0, c6288_wire_1417_0});
or_n #(2, 0, 0) OR_124 (c6288_wire_1416, {c6288_wire_1414, c6288_wire_1418});
and_n #(2, 0, 0) AND_656 (c6288_wire_1419, {c6288_wire_1416_1, c6288_wire_1417_1});
notg #(0, 0) NOT_142 (c6288_wire_1418, c6288_wire_1420);
and_n #(2, 0, 0) AND_657 (c6288_wire_1421, {c6288_wire_1422_0, c6288_wire_1423_0});
or_n #(2, 0, 0) OR_125 (c6288_wire_1422, {c6288_wire_1346, c6288_wire_1419});
and_n #(2, 0, 0) AND_658 (c6288_wire_1424, {c6288_wire_1422_1, c6288_wire_1423_1});
xor_n #(2, 0, 0) XOR_105 (c6288_wire_484, {c6288_wire_1425_0, c6288_wire_1426_0});
or_n #(2, 0, 0) OR_126 (c6288_wire_1425, {c6288_wire_1427, c6288_wire_1428});
and_n #(2, 0, 0) AND_659 (c6288_wire_1429, {c6288_wire_1425_1, c6288_wire_1426_1});
and_n #(2, 0, 0) AND_660 (c6288_wire_1428, {c6288_wire_1392, c6288_wire_1391_1});
notg #(0, 0) NOT_143 (c6288_wire_1427, c6288_wire_1430);
xor_n #(2, 0, 0) XOR_106 (c6288_wire_482, {c6288_wire_1431_0, c6288_wire_1432_0});
or_n #(2, 0, 0) OR_127 (c6288_wire_1431, {c6288_wire_1429, c6288_wire_1433});
and_n #(2, 0, 0) AND_661 (c6288_wire_1434, {c6288_wire_1431_1, c6288_wire_1432_1});
notg #(0, 0) NOT_144 (c6288_wire_1433, c6288_wire_1435);
xor_n #(2, 0, 0) XOR_107 (c6288_wire_480, {c6288_wire_1436_0, c6288_wire_1437_0});
or_n #(2, 0, 0) OR_128 (c6288_wire_1436, {c6288_wire_1434, c6288_wire_1438});
and_n #(2, 0, 0) AND_662 (c6288_wire_1439, {c6288_wire_1436_1, c6288_wire_1437_1});
notg #(0, 0) NOT_145 (c6288_wire_1438, c6288_wire_1440);
xor_n #(2, 0, 0) XOR_108 (c6288_wire_478, {c6288_wire_1441_0, c6288_wire_1442_0});
or_n #(2, 0, 0) OR_129 (c6288_wire_1441, {c6288_wire_1439, c6288_wire_1443});
and_n #(2, 0, 0) AND_663 (c6288_wire_1444, {c6288_wire_1441_1, c6288_wire_1442_1});
notg #(0, 0) NOT_146 (c6288_wire_1443, c6288_wire_1445);
xor_n #(2, 0, 0) XOR_109 (c6288_wire_476, {c6288_wire_1446_0, c6288_wire_1447_0});
or_n #(2, 0, 0) OR_130 (c6288_wire_1446, {c6288_wire_1444, c6288_wire_1448});
and_n #(2, 0, 0) AND_664 (c6288_wire_1449, {c6288_wire_1446_1, c6288_wire_1447_1});
notg #(0, 0) NOT_147 (c6288_wire_1448, c6288_wire_1450);
xor_n #(2, 0, 0) XOR_110 (c6288_wire_474, {c6288_wire_1451_0, c6288_wire_1452_0});
or_n #(2, 0, 0) OR_131 (c6288_wire_1451, {c6288_wire_1449, c6288_wire_1453});
and_n #(2, 0, 0) AND_665 (c6288_wire_1454, {c6288_wire_1451_1, c6288_wire_1452_1});
notg #(0, 0) NOT_148 (c6288_wire_1453, c6288_wire_1455);
xor_n #(2, 0, 0) XOR_111 (c6288_wire_472, {c6288_wire_1456_0, c6288_wire_1457_0});
or_n #(2, 0, 0) OR_132 (c6288_wire_1456, {c6288_wire_1454, c6288_wire_1458});
and_n #(2, 0, 0) AND_666 (c6288_wire_1459, {c6288_wire_1456_1, c6288_wire_1457_1});
notg #(0, 0) NOT_149 (c6288_wire_1458, c6288_wire_1460);
xor_n #(2, 0, 0) XOR_112 (c6288_wire_470, {c6288_wire_1461_0, c6288_wire_1462_0});
or_n #(2, 0, 0) OR_133 (c6288_wire_1461, {c6288_wire_1459, c6288_wire_1463});
and_n #(2, 0, 0) AND_667 (c6288_wire_1464, {c6288_wire_1461_1, c6288_wire_1462_1});
notg #(0, 0) NOT_150 (c6288_wire_1463, c6288_wire_1465);
xor_n #(2, 0, 0) XOR_113 (c6288_wire_468, {c6288_wire_1398_1, c6288_wire_1399_1});
or_n #(2, 0, 0) OR_134 (c6288_wire_1398, {c6288_wire_1464, c6288_wire_1466});
notg #(0, 0) NOT_151 (c6288_wire_1466, c6288_wire_1467);
and_n #(2, 0, 0) AND_668 (c6288_wire_1468, {c6288_wire_53_0, c6288_wire_1469_0});
notg #(0, 0) NOT_152 (c6288_wire_1470, c6288_wire_53_1);
xor_n #(2, 0, 0) XOR_114 (c6288_wire_508, {c6288_wire_1471_0, c6288_wire_1472_0});
or_n #(2, 0, 0) OR_135 (c6288_wire_1471, {c6288_wire_1473, c6288_wire_1474});
and_n #(2, 0, 0) AND_669 (c6288_wire_1475, {c6288_wire_1471_1, c6288_wire_1472_1});
and_n #(2, 0, 0) AND_670 (c6288_wire_1473, {c6288_wire_1476_0, c6288_wire_1477_0});
notg #(0, 0) NOT_153 (c6288_wire_1474, c6288_wire_1478);
xor_n #(2, 0, 0) XOR_115 (c6288_wire_506, {c6288_wire_1479_0, c6288_wire_1480_0});
or_n #(2, 0, 0) OR_136 (c6288_wire_1479, {c6288_wire_1475, c6288_wire_1481});
and_n #(2, 0, 0) AND_671 (c6288_wire_1482, {c6288_wire_1479_1, c6288_wire_1480_1});
notg #(0, 0) NOT_154 (c6288_wire_1481, c6288_wire_1483);
xor_n #(2, 0, 0) XOR_116 (c6288_wire_504, {c6288_wire_1484_0, c6288_wire_1485_0});
or_n #(2, 0, 0) OR_137 (c6288_wire_1484, {c6288_wire_1482, c6288_wire_1486});
and_n #(2, 0, 0) AND_672 (c6288_wire_1487, {c6288_wire_1484_1, c6288_wire_1485_1});
notg #(0, 0) NOT_155 (c6288_wire_1486, c6288_wire_1488);
xor_n #(2, 0, 0) XOR_117 (c6288_wire_502, {c6288_wire_1489_0, c6288_wire_1490_0});
or_n #(2, 0, 0) OR_138 (c6288_wire_1489, {c6288_wire_1487, c6288_wire_1491});
and_n #(2, 0, 0) AND_673 (c6288_wire_1492, {c6288_wire_1489_1, c6288_wire_1490_1});
notg #(0, 0) NOT_156 (c6288_wire_1491, c6288_wire_1493);
xor_n #(2, 0, 0) XOR_118 (c6288_wire_1423, {c6288_wire_1494_0, c6288_wire_1495_0});
or_n #(2, 0, 0) OR_139 (c6288_wire_1494, {c6288_wire_1492, c6288_wire_1496});
and_n #(2, 0, 0) AND_674 (c6288_wire_1497, {c6288_wire_1494_1, c6288_wire_1495_1});
notg #(0, 0) NOT_157 (c6288_wire_1496, c6288_wire_1498);
and_n #(2, 0, 0) AND_675 (c6288_wire_1499, {c6288_wire_1500_0, c6288_wire_1501_0});
or_n #(2, 0, 0) OR_140 (c6288_wire_1500, {c6288_wire_1424, c6288_wire_1497});
and_n #(2, 0, 0) AND_676 (c6288_wire_1502, {c6288_wire_1500_1, c6288_wire_1501_1});
xor_n #(2, 0, 0) XOR_119 (c6288_wire_526, {c6288_wire_1503_0, c6288_wire_1504_0});
or_n #(2, 0, 0) OR_141 (c6288_wire_1503, {c6288_wire_1505, c6288_wire_1506});
and_n #(2, 0, 0) AND_677 (c6288_wire_1507, {c6288_wire_1503_1, c6288_wire_1504_1});
and_n #(2, 0, 0) AND_678 (c6288_wire_1506, {c6288_wire_1470, c6288_wire_1469_1});
notg #(0, 0) NOT_158 (c6288_wire_1505, c6288_wire_1508);
xor_n #(2, 0, 0) XOR_120 (c6288_wire_524, {c6288_wire_1509_0, c6288_wire_1510_0});
or_n #(2, 0, 0) OR_142 (c6288_wire_1509, {c6288_wire_1507, c6288_wire_1511});
and_n #(2, 0, 0) AND_679 (c6288_wire_1512, {c6288_wire_1509_1, c6288_wire_1510_1});
notg #(0, 0) NOT_159 (c6288_wire_1511, c6288_wire_1513);
xor_n #(2, 0, 0) XOR_121 (c6288_wire_522, {c6288_wire_1514_0, c6288_wire_1515_0});
or_n #(2, 0, 0) OR_143 (c6288_wire_1514, {c6288_wire_1512, c6288_wire_1516});
and_n #(2, 0, 0) AND_680 (c6288_wire_1517, {c6288_wire_1514_1, c6288_wire_1515_1});
notg #(0, 0) NOT_160 (c6288_wire_1516, c6288_wire_1518);
xor_n #(2, 0, 0) XOR_122 (c6288_wire_520, {c6288_wire_1519_0, c6288_wire_1520_0});
or_n #(2, 0, 0) OR_144 (c6288_wire_1519, {c6288_wire_1517, c6288_wire_1521});
and_n #(2, 0, 0) AND_681 (c6288_wire_1522, {c6288_wire_1519_1, c6288_wire_1520_1});
notg #(0, 0) NOT_161 (c6288_wire_1521, c6288_wire_1523);
xor_n #(2, 0, 0) XOR_123 (c6288_wire_518, {c6288_wire_1524_0, c6288_wire_1525_0});
or_n #(2, 0, 0) OR_145 (c6288_wire_1524, {c6288_wire_1522, c6288_wire_1526});
and_n #(2, 0, 0) AND_682 (c6288_wire_1527, {c6288_wire_1524_1, c6288_wire_1525_1});
notg #(0, 0) NOT_162 (c6288_wire_1526, c6288_wire_1528);
xor_n #(2, 0, 0) XOR_124 (c6288_wire_516, {c6288_wire_1529_0, c6288_wire_1530_0});
or_n #(2, 0, 0) OR_146 (c6288_wire_1529, {c6288_wire_1527, c6288_wire_1531});
and_n #(2, 0, 0) AND_683 (c6288_wire_1532, {c6288_wire_1529_1, c6288_wire_1530_1});
notg #(0, 0) NOT_163 (c6288_wire_1531, c6288_wire_1533);
xor_n #(2, 0, 0) XOR_125 (c6288_wire_514, {c6288_wire_1534_0, c6288_wire_1535_0});
or_n #(2, 0, 0) OR_147 (c6288_wire_1534, {c6288_wire_1532, c6288_wire_1536});
and_n #(2, 0, 0) AND_684 (c6288_wire_1537, {c6288_wire_1534_1, c6288_wire_1535_1});
notg #(0, 0) NOT_164 (c6288_wire_1536, c6288_wire_1538);
xor_n #(2, 0, 0) XOR_126 (c6288_wire_512, {c6288_wire_1539_0, c6288_wire_1540_0});
or_n #(2, 0, 0) OR_148 (c6288_wire_1539, {c6288_wire_1537, c6288_wire_1541});
and_n #(2, 0, 0) AND_685 (c6288_wire_1542, {c6288_wire_1539_1, c6288_wire_1540_1});
notg #(0, 0) NOT_165 (c6288_wire_1541, c6288_wire_1543);
xor_n #(2, 0, 0) XOR_127 (c6288_wire_510, {c6288_wire_1476_1, c6288_wire_1477_1});
or_n #(2, 0, 0) OR_149 (c6288_wire_1476, {c6288_wire_1542, c6288_wire_1544});
notg #(0, 0) NOT_166 (c6288_wire_1544, c6288_wire_1545);
and_n #(2, 0, 0) AND_686 (c6288_wire_1546, {c6288_wire_58_0, c6288_wire_1547_0});
notg #(0, 0) NOT_167 (c6288_wire_1548, c6288_wire_58_1);
xor_n #(2, 0, 0) XOR_128 (c6288_wire_550, {c6288_wire_1549_0, c6288_wire_1550_0});
or_n #(2, 0, 0) OR_150 (c6288_wire_1549, {c6288_wire_1551, c6288_wire_1552});
and_n #(2, 0, 0) AND_687 (c6288_wire_1553, {c6288_wire_1549_1, c6288_wire_1550_1});
and_n #(2, 0, 0) AND_688 (c6288_wire_1551, {c6288_wire_1554_0, c6288_wire_1555_0});
notg #(0, 0) NOT_168 (c6288_wire_1552, c6288_wire_1556);
xor_n #(2, 0, 0) XOR_129 (c6288_wire_548, {c6288_wire_1557_0, c6288_wire_1558_0});
or_n #(2, 0, 0) OR_151 (c6288_wire_1557, {c6288_wire_1553, c6288_wire_1559});
and_n #(2, 0, 0) AND_689 (c6288_wire_1560, {c6288_wire_1557_1, c6288_wire_1558_1});
notg #(0, 0) NOT_169 (c6288_wire_1559, c6288_wire_1561);
xor_n #(2, 0, 0) XOR_130 (c6288_wire_546, {c6288_wire_1562_0, c6288_wire_1563_0});
or_n #(2, 0, 0) OR_152 (c6288_wire_1562, {c6288_wire_1560, c6288_wire_1564});
and_n #(2, 0, 0) AND_690 (c6288_wire_1565, {c6288_wire_1562_1, c6288_wire_1563_1});
notg #(0, 0) NOT_170 (c6288_wire_1564, c6288_wire_1566);
xor_n #(2, 0, 0) XOR_131 (c6288_wire_544, {c6288_wire_1567_0, c6288_wire_1568_0});
or_n #(2, 0, 0) OR_153 (c6288_wire_1567, {c6288_wire_1565, c6288_wire_1569});
and_n #(2, 0, 0) AND_691 (c6288_wire_1570, {c6288_wire_1567_1, c6288_wire_1568_1});
notg #(0, 0) NOT_171 (c6288_wire_1569, c6288_wire_1571);
xor_n #(2, 0, 0) XOR_132 (c6288_wire_1501, {c6288_wire_1572_0, c6288_wire_1573_0});
or_n #(2, 0, 0) OR_154 (c6288_wire_1572, {c6288_wire_1570, c6288_wire_1574});
and_n #(2, 0, 0) AND_692 (c6288_wire_1575, {c6288_wire_1572_1, c6288_wire_1573_1});
notg #(0, 0) NOT_172 (c6288_wire_1574, c6288_wire_1576);
and_n #(2, 0, 0) AND_693 (c6288_wire_1577, {c6288_wire_1578_0, c6288_wire_1579_0});
or_n #(2, 0, 0) OR_155 (c6288_wire_1578, {c6288_wire_1502, c6288_wire_1575});
and_n #(2, 0, 0) AND_694 (c6288_wire_1580, {c6288_wire_1578_1, c6288_wire_1579_1});
xor_n #(2, 0, 0) XOR_133 (c6288_wire_568, {c6288_wire_1581_0, c6288_wire_1582_0});
or_n #(2, 0, 0) OR_156 (c6288_wire_1581, {c6288_wire_1583, c6288_wire_1584});
and_n #(2, 0, 0) AND_695 (c6288_wire_1585, {c6288_wire_1581_1, c6288_wire_1582_1});
and_n #(2, 0, 0) AND_696 (c6288_wire_1584, {c6288_wire_1548, c6288_wire_1547_1});
notg #(0, 0) NOT_173 (c6288_wire_1583, c6288_wire_1586);
xor_n #(2, 0, 0) XOR_134 (c6288_wire_566, {c6288_wire_1587_0, c6288_wire_1588_0});
or_n #(2, 0, 0) OR_157 (c6288_wire_1587, {c6288_wire_1585, c6288_wire_1589});
and_n #(2, 0, 0) AND_697 (c6288_wire_1590, {c6288_wire_1587_1, c6288_wire_1588_1});
notg #(0, 0) NOT_174 (c6288_wire_1589, c6288_wire_1591);
xor_n #(2, 0, 0) XOR_135 (c6288_wire_564, {c6288_wire_1592_0, c6288_wire_1593_0});
or_n #(2, 0, 0) OR_158 (c6288_wire_1592, {c6288_wire_1590, c6288_wire_1594});
and_n #(2, 0, 0) AND_698 (c6288_wire_1595, {c6288_wire_1592_1, c6288_wire_1593_1});
notg #(0, 0) NOT_175 (c6288_wire_1594, c6288_wire_1596);
xor_n #(2, 0, 0) XOR_136 (c6288_wire_562, {c6288_wire_1597_0, c6288_wire_1598_0});
or_n #(2, 0, 0) OR_159 (c6288_wire_1597, {c6288_wire_1595, c6288_wire_1599});
and_n #(2, 0, 0) AND_699 (c6288_wire_1600, {c6288_wire_1597_1, c6288_wire_1598_1});
notg #(0, 0) NOT_176 (c6288_wire_1599, c6288_wire_1601);
xor_n #(2, 0, 0) XOR_137 (c6288_wire_560, {c6288_wire_1602_0, c6288_wire_1603_0});
or_n #(2, 0, 0) OR_160 (c6288_wire_1602, {c6288_wire_1600, c6288_wire_1604});
and_n #(2, 0, 0) AND_700 (c6288_wire_1605, {c6288_wire_1602_1, c6288_wire_1603_1});
notg #(0, 0) NOT_177 (c6288_wire_1604, c6288_wire_1606);
xor_n #(2, 0, 0) XOR_138 (c6288_wire_558, {c6288_wire_1607_0, c6288_wire_1608_0});
or_n #(2, 0, 0) OR_161 (c6288_wire_1607, {c6288_wire_1605, c6288_wire_1609});
and_n #(2, 0, 0) AND_701 (c6288_wire_1610, {c6288_wire_1607_1, c6288_wire_1608_1});
notg #(0, 0) NOT_178 (c6288_wire_1609, c6288_wire_1611);
xor_n #(2, 0, 0) XOR_139 (c6288_wire_556, {c6288_wire_1612_0, c6288_wire_1613_0});
or_n #(2, 0, 0) OR_162 (c6288_wire_1612, {c6288_wire_1610, c6288_wire_1614});
and_n #(2, 0, 0) AND_702 (c6288_wire_1615, {c6288_wire_1612_1, c6288_wire_1613_1});
notg #(0, 0) NOT_179 (c6288_wire_1614, c6288_wire_1616);
xor_n #(2, 0, 0) XOR_140 (c6288_wire_554, {c6288_wire_1617_0, c6288_wire_1618_0});
or_n #(2, 0, 0) OR_163 (c6288_wire_1617, {c6288_wire_1615, c6288_wire_1619});
and_n #(2, 0, 0) AND_703 (c6288_wire_1620, {c6288_wire_1617_1, c6288_wire_1618_1});
notg #(0, 0) NOT_180 (c6288_wire_1619, c6288_wire_1621);
xor_n #(2, 0, 0) XOR_141 (c6288_wire_552, {c6288_wire_1554_1, c6288_wire_1555_1});
or_n #(2, 0, 0) OR_164 (c6288_wire_1554, {c6288_wire_1620, c6288_wire_1622});
notg #(0, 0) NOT_181 (c6288_wire_1622, c6288_wire_1623);
and_n #(2, 0, 0) AND_704 (c6288_wire_1624, {c6288_wire_63_0, c6288_wire_1625_0});
notg #(0, 0) NOT_182 (c6288_wire_1626, c6288_wire_63_1);
xor_n #(2, 0, 0) XOR_142 (c6288_wire_592, {c6288_wire_1627_0, c6288_wire_1628_0});
or_n #(2, 0, 0) OR_165 (c6288_wire_1627, {c6288_wire_1629, c6288_wire_1630});
and_n #(2, 0, 0) AND_705 (c6288_wire_1631, {c6288_wire_1627_1, c6288_wire_1628_1});
and_n #(2, 0, 0) AND_706 (c6288_wire_1629, {c6288_wire_1632_0, c6288_wire_1633_0});
notg #(0, 0) NOT_183 (c6288_wire_1630, c6288_wire_1634);
xor_n #(2, 0, 0) XOR_143 (c6288_wire_590, {c6288_wire_1635_0, c6288_wire_1636_0});
or_n #(2, 0, 0) OR_166 (c6288_wire_1635, {c6288_wire_1631, c6288_wire_1637});
and_n #(2, 0, 0) AND_707 (c6288_wire_1638, {c6288_wire_1635_1, c6288_wire_1636_1});
notg #(0, 0) NOT_184 (c6288_wire_1637, c6288_wire_1639);
xor_n #(2, 0, 0) XOR_144 (c6288_wire_588, {c6288_wire_1640_0, c6288_wire_1641_0});
or_n #(2, 0, 0) OR_167 (c6288_wire_1640, {c6288_wire_1638, c6288_wire_1642});
and_n #(2, 0, 0) AND_708 (c6288_wire_1643, {c6288_wire_1640_1, c6288_wire_1641_1});
notg #(0, 0) NOT_185 (c6288_wire_1642, c6288_wire_1644);
xor_n #(2, 0, 0) XOR_145 (c6288_wire_586, {c6288_wire_1645_0, c6288_wire_1646_0});
or_n #(2, 0, 0) OR_168 (c6288_wire_1645, {c6288_wire_1643, c6288_wire_1647});
and_n #(2, 0, 0) AND_709 (c6288_wire_1648, {c6288_wire_1645_1, c6288_wire_1646_1});
notg #(0, 0) NOT_186 (c6288_wire_1647, c6288_wire_1649);
xor_n #(2, 0, 0) XOR_146 (c6288_wire_1579, {c6288_wire_1650_0, c6288_wire_1651_0});
or_n #(2, 0, 0) OR_169 (c6288_wire_1650, {c6288_wire_1648, c6288_wire_1652});
and_n #(2, 0, 0) AND_710 (c6288_wire_1653, {c6288_wire_1650_1, c6288_wire_1651_1});
notg #(0, 0) NOT_187 (c6288_wire_1652, c6288_wire_1654);
and_n #(2, 0, 0) AND_711 (c6288_wire_1655, {c6288_wire_1656_0, c6288_wire_1657_0});
or_n #(2, 0, 0) OR_170 (c6288_wire_1656, {c6288_wire_1580, c6288_wire_1653});
and_n #(2, 0, 0) AND_712 (c6288_wire_1658, {c6288_wire_1656_1, c6288_wire_1657_1});
xor_n #(2, 0, 0) XOR_147 (c6288_wire_610, {c6288_wire_1659_0, c6288_wire_1660_0});
or_n #(2, 0, 0) OR_171 (c6288_wire_1659, {c6288_wire_1661, c6288_wire_1662});
and_n #(2, 0, 0) AND_713 (c6288_wire_1663, {c6288_wire_1659_1, c6288_wire_1660_1});
and_n #(2, 0, 0) AND_714 (c6288_wire_1662, {c6288_wire_1626, c6288_wire_1625_1});
notg #(0, 0) NOT_188 (c6288_wire_1661, c6288_wire_1664);
xor_n #(2, 0, 0) XOR_148 (c6288_wire_608, {c6288_wire_1665_0, c6288_wire_1666_0});
or_n #(2, 0, 0) OR_172 (c6288_wire_1665, {c6288_wire_1663, c6288_wire_1667});
and_n #(2, 0, 0) AND_715 (c6288_wire_1668, {c6288_wire_1665_1, c6288_wire_1666_1});
notg #(0, 0) NOT_189 (c6288_wire_1667, c6288_wire_1669);
xor_n #(2, 0, 0) XOR_149 (c6288_wire_606, {c6288_wire_1670_0, c6288_wire_1671_0});
or_n #(2, 0, 0) OR_173 (c6288_wire_1670, {c6288_wire_1668, c6288_wire_1672});
and_n #(2, 0, 0) AND_716 (c6288_wire_1673, {c6288_wire_1670_1, c6288_wire_1671_1});
notg #(0, 0) NOT_190 (c6288_wire_1672, c6288_wire_1674);
xor_n #(2, 0, 0) XOR_150 (c6288_wire_604, {c6288_wire_1675_0, c6288_wire_1676_0});
or_n #(2, 0, 0) OR_174 (c6288_wire_1675, {c6288_wire_1673, c6288_wire_1677});
and_n #(2, 0, 0) AND_717 (c6288_wire_1678, {c6288_wire_1675_1, c6288_wire_1676_1});
notg #(0, 0) NOT_191 (c6288_wire_1677, c6288_wire_1679);
xor_n #(2, 0, 0) XOR_151 (c6288_wire_602, {c6288_wire_1680_0, c6288_wire_1681_0});
or_n #(2, 0, 0) OR_175 (c6288_wire_1680, {c6288_wire_1678, c6288_wire_1682});
and_n #(2, 0, 0) AND_718 (c6288_wire_1683, {c6288_wire_1680_1, c6288_wire_1681_1});
notg #(0, 0) NOT_192 (c6288_wire_1682, c6288_wire_1684);
xor_n #(2, 0, 0) XOR_152 (c6288_wire_600, {c6288_wire_1685_0, c6288_wire_1686_0});
or_n #(2, 0, 0) OR_176 (c6288_wire_1685, {c6288_wire_1683, c6288_wire_1687});
and_n #(2, 0, 0) AND_719 (c6288_wire_1688, {c6288_wire_1685_1, c6288_wire_1686_1});
notg #(0, 0) NOT_193 (c6288_wire_1687, c6288_wire_1689);
xor_n #(2, 0, 0) XOR_153 (c6288_wire_598, {c6288_wire_1690_0, c6288_wire_1691_0});
or_n #(2, 0, 0) OR_177 (c6288_wire_1690, {c6288_wire_1688, c6288_wire_1692});
and_n #(2, 0, 0) AND_720 (c6288_wire_1693, {c6288_wire_1690_1, c6288_wire_1691_1});
notg #(0, 0) NOT_194 (c6288_wire_1692, c6288_wire_1694);
xor_n #(2, 0, 0) XOR_154 (c6288_wire_596, {c6288_wire_1695_0, c6288_wire_1696_0});
or_n #(2, 0, 0) OR_178 (c6288_wire_1695, {c6288_wire_1693, c6288_wire_1697});
and_n #(2, 0, 0) AND_721 (c6288_wire_1698, {c6288_wire_1695_1, c6288_wire_1696_1});
notg #(0, 0) NOT_195 (c6288_wire_1697, c6288_wire_1699);
xor_n #(2, 0, 0) XOR_155 (c6288_wire_594, {c6288_wire_1632_1, c6288_wire_1633_1});
or_n #(2, 0, 0) OR_179 (c6288_wire_1632, {c6288_wire_1698, c6288_wire_1700});
notg #(0, 0) NOT_196 (c6288_wire_1700, c6288_wire_1701);
and_n #(2, 0, 0) AND_722 (c6288_wire_1702, {c6288_wire_68_0, c6288_wire_1703_0});
notg #(0, 0) NOT_197 (c6288_wire_1704, c6288_wire_68_1);
xor_n #(2, 0, 0) XOR_156 (c6288_wire_634, {c6288_wire_1705_0, c6288_wire_1706_0});
or_n #(2, 0, 0) OR_180 (c6288_wire_1705, {c6288_wire_1707, c6288_wire_1708});
and_n #(2, 0, 0) AND_723 (c6288_wire_1709, {c6288_wire_1705_1, c6288_wire_1706_1});
and_n #(2, 0, 0) AND_724 (c6288_wire_1707, {c6288_wire_1710_0, c6288_wire_1711_0});
notg #(0, 0) NOT_198 (c6288_wire_1708, c6288_wire_1712);
xor_n #(2, 0, 0) XOR_157 (c6288_wire_632, {c6288_wire_1713_0, c6288_wire_1714_0});
or_n #(2, 0, 0) OR_181 (c6288_wire_1713, {c6288_wire_1709, c6288_wire_1715});
and_n #(2, 0, 0) AND_725 (c6288_wire_1716, {c6288_wire_1713_1, c6288_wire_1714_1});
notg #(0, 0) NOT_199 (c6288_wire_1715, c6288_wire_1717);
xor_n #(2, 0, 0) XOR_158 (c6288_wire_630, {c6288_wire_1718_0, c6288_wire_1719_0});
or_n #(2, 0, 0) OR_182 (c6288_wire_1718, {c6288_wire_1716, c6288_wire_1720});
and_n #(2, 0, 0) AND_726 (c6288_wire_1721, {c6288_wire_1718_1, c6288_wire_1719_1});
notg #(0, 0) NOT_200 (c6288_wire_1720, c6288_wire_1722);
xor_n #(2, 0, 0) XOR_159 (c6288_wire_628, {c6288_wire_1723_0, c6288_wire_1724_0});
or_n #(2, 0, 0) OR_183 (c6288_wire_1723, {c6288_wire_1721, c6288_wire_1725});
and_n #(2, 0, 0) AND_727 (c6288_wire_1726, {c6288_wire_1723_1, c6288_wire_1724_1});
notg #(0, 0) NOT_201 (c6288_wire_1725, c6288_wire_1727);
xor_n #(2, 0, 0) XOR_160 (c6288_wire_1657, {c6288_wire_1728_0, c6288_wire_1729_0});
or_n #(2, 0, 0) OR_184 (c6288_wire_1728, {c6288_wire_1726, c6288_wire_1730});
and_n #(2, 0, 0) AND_728 (c6288_wire_1731, {c6288_wire_1728_1, c6288_wire_1729_1});
notg #(0, 0) NOT_202 (c6288_wire_1730, c6288_wire_1732);
and_n #(2, 0, 0) AND_729 (c6288_wire_1733, {c6288_wire_1734_0, c6288_wire_1735_0});
or_n #(2, 0, 0) OR_185 (c6288_wire_1734, {c6288_wire_1658, c6288_wire_1731});
and_n #(2, 0, 0) AND_730 (c6288_wire_1736, {c6288_wire_1734_1, c6288_wire_1735_1});
xor_n #(2, 0, 0) XOR_161 (c6288_wire_652, {c6288_wire_1737_0, c6288_wire_1738_0});
or_n #(2, 0, 0) OR_186 (c6288_wire_1737, {c6288_wire_1739, c6288_wire_1740});
and_n #(2, 0, 0) AND_731 (c6288_wire_1741, {c6288_wire_1737_1, c6288_wire_1738_1});
and_n #(2, 0, 0) AND_732 (c6288_wire_1740, {c6288_wire_1704, c6288_wire_1703_1});
notg #(0, 0) NOT_203 (c6288_wire_1739, c6288_wire_1742);
xor_n #(2, 0, 0) XOR_162 (c6288_wire_650, {c6288_wire_1743_0, c6288_wire_1744_0});
or_n #(2, 0, 0) OR_187 (c6288_wire_1743, {c6288_wire_1741, c6288_wire_1745});
and_n #(2, 0, 0) AND_733 (c6288_wire_1746, {c6288_wire_1743_1, c6288_wire_1744_1});
notg #(0, 0) NOT_204 (c6288_wire_1745, c6288_wire_1747);
xor_n #(2, 0, 0) XOR_163 (c6288_wire_648, {c6288_wire_1748_0, c6288_wire_1749_0});
or_n #(2, 0, 0) OR_188 (c6288_wire_1748, {c6288_wire_1746, c6288_wire_1750});
and_n #(2, 0, 0) AND_734 (c6288_wire_1751, {c6288_wire_1748_1, c6288_wire_1749_1});
notg #(0, 0) NOT_205 (c6288_wire_1750, c6288_wire_1752);
xor_n #(2, 0, 0) XOR_164 (c6288_wire_646, {c6288_wire_1753_0, c6288_wire_1754_0});
or_n #(2, 0, 0) OR_189 (c6288_wire_1753, {c6288_wire_1751, c6288_wire_1755});
and_n #(2, 0, 0) AND_735 (c6288_wire_1756, {c6288_wire_1753_1, c6288_wire_1754_1});
notg #(0, 0) NOT_206 (c6288_wire_1755, c6288_wire_1757);
xor_n #(2, 0, 0) XOR_165 (c6288_wire_644, {c6288_wire_1758_0, c6288_wire_1759_0});
or_n #(2, 0, 0) OR_190 (c6288_wire_1758, {c6288_wire_1756, c6288_wire_1760});
and_n #(2, 0, 0) AND_736 (c6288_wire_1761, {c6288_wire_1758_1, c6288_wire_1759_1});
notg #(0, 0) NOT_207 (c6288_wire_1760, c6288_wire_1762);
xor_n #(2, 0, 0) XOR_166 (c6288_wire_642, {c6288_wire_1763_0, c6288_wire_1764_0});
or_n #(2, 0, 0) OR_191 (c6288_wire_1763, {c6288_wire_1761, c6288_wire_1765});
and_n #(2, 0, 0) AND_737 (c6288_wire_1766, {c6288_wire_1763_1, c6288_wire_1764_1});
notg #(0, 0) NOT_208 (c6288_wire_1765, c6288_wire_1767);
xor_n #(2, 0, 0) XOR_167 (c6288_wire_640, {c6288_wire_1768_0, c6288_wire_1769_0});
or_n #(2, 0, 0) OR_192 (c6288_wire_1768, {c6288_wire_1766, c6288_wire_1770});
and_n #(2, 0, 0) AND_738 (c6288_wire_1771, {c6288_wire_1768_1, c6288_wire_1769_1});
notg #(0, 0) NOT_209 (c6288_wire_1770, c6288_wire_1772);
xor_n #(2, 0, 0) XOR_168 (c6288_wire_638, {c6288_wire_1773_0, c6288_wire_1774_0});
or_n #(2, 0, 0) OR_193 (c6288_wire_1773, {c6288_wire_1771, c6288_wire_1775});
and_n #(2, 0, 0) AND_739 (c6288_wire_1776, {c6288_wire_1773_1, c6288_wire_1774_1});
notg #(0, 0) NOT_210 (c6288_wire_1775, c6288_wire_1777);
xor_n #(2, 0, 0) XOR_169 (c6288_wire_636, {c6288_wire_1710_1, c6288_wire_1711_1});
or_n #(2, 0, 0) OR_194 (c6288_wire_1710, {c6288_wire_1776, c6288_wire_1778});
notg #(0, 0) NOT_211 (c6288_wire_1778, c6288_wire_1779);
and_n #(2, 0, 0) AND_740 (c6288_wire_1780, {c6288_wire_72_0, c6288_wire_1781_0});
notg #(0, 0) NOT_212 (c6288_wire_1782, c6288_wire_72_1);
xor_n #(2, 0, 0) XOR_170 (c6288_wire_676, {c6288_wire_1783_0, c6288_wire_1784_0});
or_n #(2, 0, 0) OR_195 (c6288_wire_1783, {c6288_wire_1785, c6288_wire_1786});
and_n #(2, 0, 0) AND_741 (c6288_wire_1787, {c6288_wire_1783_1, c6288_wire_1784_1});
and_n #(2, 0, 0) AND_742 (c6288_wire_1785, {c6288_wire_1788_0, c6288_wire_1789_0});
notg #(0, 0) NOT_213 (c6288_wire_1786, c6288_wire_1790);
xor_n #(2, 0, 0) XOR_171 (c6288_wire_674, {c6288_wire_1791_0, c6288_wire_1792_0});
or_n #(2, 0, 0) OR_196 (c6288_wire_1791, {c6288_wire_1787, c6288_wire_1793});
and_n #(2, 0, 0) AND_743 (c6288_wire_1794, {c6288_wire_1791_1, c6288_wire_1792_1});
notg #(0, 0) NOT_214 (c6288_wire_1793, c6288_wire_1795);
xor_n #(2, 0, 0) XOR_172 (c6288_wire_672, {c6288_wire_1796_0, c6288_wire_1797_0});
or_n #(2, 0, 0) OR_197 (c6288_wire_1796, {c6288_wire_1794, c6288_wire_1798});
and_n #(2, 0, 0) AND_744 (c6288_wire_1799, {c6288_wire_1796_1, c6288_wire_1797_1});
notg #(0, 0) NOT_215 (c6288_wire_1798, c6288_wire_1800);
xor_n #(2, 0, 0) XOR_173 (c6288_wire_670, {c6288_wire_1801_0, c6288_wire_1802_0});
or_n #(2, 0, 0) OR_198 (c6288_wire_1801, {c6288_wire_1799, c6288_wire_1803});
and_n #(2, 0, 0) AND_745 (c6288_wire_1804, {c6288_wire_1801_1, c6288_wire_1802_1});
notg #(0, 0) NOT_216 (c6288_wire_1803, c6288_wire_1805);
xor_n #(2, 0, 0) XOR_174 (c6288_wire_1735, {c6288_wire_1806_0, c6288_wire_1807_0});
or_n #(2, 0, 0) OR_199 (c6288_wire_1806, {c6288_wire_1804, c6288_wire_1808});
and_n #(2, 0, 0) AND_746 (c6288_wire_1809, {c6288_wire_1806_1, c6288_wire_1807_1});
notg #(0, 0) NOT_217 (c6288_wire_1808, c6288_wire_1810);
and_n #(2, 0, 0) AND_747 (c6288_wire_1811, {c6288_wire_1812_0, c6288_wire_1813_0});
or_n #(2, 0, 0) OR_200 (c6288_wire_1812, {c6288_wire_1736, c6288_wire_1809});
and_n #(2, 0, 0) AND_748 (c6288_wire_1814, {c6288_wire_1812_1, c6288_wire_1813_1});
xor_n #(2, 0, 0) XOR_175 (c6288_wire_694, {c6288_wire_1815_0, c6288_wire_1816_0});
or_n #(2, 0, 0) OR_201 (c6288_wire_1815, {c6288_wire_1817, c6288_wire_1818});
and_n #(2, 0, 0) AND_749 (c6288_wire_1819, {c6288_wire_1815_1, c6288_wire_1816_1});
and_n #(2, 0, 0) AND_750 (c6288_wire_1818, {c6288_wire_1782, c6288_wire_1781_1});
notg #(0, 0) NOT_218 (c6288_wire_1817, c6288_wire_1820);
xor_n #(2, 0, 0) XOR_176 (c6288_wire_692, {c6288_wire_1821_0, c6288_wire_1822_0});
or_n #(2, 0, 0) OR_202 (c6288_wire_1821, {c6288_wire_1819, c6288_wire_1823});
and_n #(2, 0, 0) AND_751 (c6288_wire_1824, {c6288_wire_1821_1, c6288_wire_1822_1});
notg #(0, 0) NOT_219 (c6288_wire_1823, c6288_wire_1825);
xor_n #(2, 0, 0) XOR_177 (c6288_wire_690, {c6288_wire_1826_0, c6288_wire_1827_0});
or_n #(2, 0, 0) OR_203 (c6288_wire_1826, {c6288_wire_1824, c6288_wire_1828});
and_n #(2, 0, 0) AND_752 (c6288_wire_1829, {c6288_wire_1826_1, c6288_wire_1827_1});
notg #(0, 0) NOT_220 (c6288_wire_1828, c6288_wire_1830);
xor_n #(2, 0, 0) XOR_178 (c6288_wire_688, {c6288_wire_1831_0, c6288_wire_1832_0});
or_n #(2, 0, 0) OR_204 (c6288_wire_1831, {c6288_wire_1829, c6288_wire_1833});
and_n #(2, 0, 0) AND_753 (c6288_wire_1834, {c6288_wire_1831_1, c6288_wire_1832_1});
notg #(0, 0) NOT_221 (c6288_wire_1833, c6288_wire_1835);
xor_n #(2, 0, 0) XOR_179 (c6288_wire_686, {c6288_wire_1836_0, c6288_wire_1837_0});
or_n #(2, 0, 0) OR_205 (c6288_wire_1836, {c6288_wire_1834, c6288_wire_1838});
and_n #(2, 0, 0) AND_754 (c6288_wire_1839, {c6288_wire_1836_1, c6288_wire_1837_1});
notg #(0, 0) NOT_222 (c6288_wire_1838, c6288_wire_1840);
xor_n #(2, 0, 0) XOR_180 (c6288_wire_684, {c6288_wire_1841_0, c6288_wire_1842_0});
or_n #(2, 0, 0) OR_206 (c6288_wire_1841, {c6288_wire_1839, c6288_wire_1843});
and_n #(2, 0, 0) AND_755 (c6288_wire_1844, {c6288_wire_1841_1, c6288_wire_1842_1});
notg #(0, 0) NOT_223 (c6288_wire_1843, c6288_wire_1845);
xor_n #(2, 0, 0) XOR_181 (c6288_wire_682, {c6288_wire_1846_0, c6288_wire_1847_0});
or_n #(2, 0, 0) OR_207 (c6288_wire_1846, {c6288_wire_1844, c6288_wire_1848});
and_n #(2, 0, 0) AND_756 (c6288_wire_1849, {c6288_wire_1846_1, c6288_wire_1847_1});
notg #(0, 0) NOT_224 (c6288_wire_1848, c6288_wire_1850);
xor_n #(2, 0, 0) XOR_182 (c6288_wire_680, {c6288_wire_1851_0, c6288_wire_1852_0});
or_n #(2, 0, 0) OR_208 (c6288_wire_1851, {c6288_wire_1849, c6288_wire_1853});
and_n #(2, 0, 0) AND_757 (c6288_wire_1854, {c6288_wire_1851_1, c6288_wire_1852_1});
notg #(0, 0) NOT_225 (c6288_wire_1853, c6288_wire_1855);
xor_n #(2, 0, 0) XOR_183 (c6288_wire_678, {c6288_wire_1788_1, c6288_wire_1789_1});
or_n #(2, 0, 0) OR_209 (c6288_wire_1788, {c6288_wire_1854, c6288_wire_1856});
notg #(0, 0) NOT_226 (c6288_wire_1856, c6288_wire_1857);
and_n #(2, 0, 0) AND_758 (c6288_wire_1858, {c6288_wire_4_0, c6288_wire_1859_0});
notg #(0, 0) NOT_227 (c6288_wire_1860, c6288_wire_4_1);
xor_n #(2, 0, 0) XOR_184 (c6288_wire_718, {c6288_wire_1861_0, c6288_wire_1862_0});
or_n #(2, 0, 0) OR_210 (c6288_wire_1861, {c6288_wire_1863, c6288_wire_1864});
and_n #(2, 0, 0) AND_759 (c6288_wire_1865, {c6288_wire_1861_1, c6288_wire_1862_1});
and_n #(2, 0, 0) AND_760 (c6288_wire_1863, {c6288_wire_1866_0, c6288_wire_1867_0});
notg #(0, 0) NOT_228 (c6288_wire_1864, c6288_wire_1868);
xor_n #(2, 0, 0) XOR_185 (c6288_wire_716, {c6288_wire_1869_0, c6288_wire_1870_0});
or_n #(2, 0, 0) OR_211 (c6288_wire_1869, {c6288_wire_1865, c6288_wire_1871});
and_n #(2, 0, 0) AND_761 (c6288_wire_1872, {c6288_wire_1869_1, c6288_wire_1870_1});
notg #(0, 0) NOT_229 (c6288_wire_1871, c6288_wire_1873);
xor_n #(2, 0, 0) XOR_186 (c6288_wire_714, {c6288_wire_1874_0, c6288_wire_1875_0});
or_n #(2, 0, 0) OR_212 (c6288_wire_1874, {c6288_wire_1872, c6288_wire_1876});
and_n #(2, 0, 0) AND_762 (c6288_wire_1877, {c6288_wire_1874_1, c6288_wire_1875_1});
notg #(0, 0) NOT_230 (c6288_wire_1876, c6288_wire_1878);
xor_n #(2, 0, 0) XOR_187 (c6288_wire_712, {c6288_wire_1879_0, c6288_wire_1880_0});
or_n #(2, 0, 0) OR_213 (c6288_wire_1879, {c6288_wire_1877, c6288_wire_1881});
and_n #(2, 0, 0) AND_763 (c6288_wire_1882, {c6288_wire_1879_1, c6288_wire_1880_1});
notg #(0, 0) NOT_231 (c6288_wire_1881, c6288_wire_1883);
xor_n #(2, 0, 0) XOR_188 (c6288_wire_1813, {c6288_wire_1884_0, c6288_wire_1885_0});
or_n #(2, 0, 0) OR_214 (c6288_wire_1884, {c6288_wire_1882, c6288_wire_1886});
and_n #(2, 0, 0) AND_764 (c6288_wire_1887, {c6288_wire_1884_1, c6288_wire_1885_1});
notg #(0, 0) NOT_232 (c6288_wire_1886, c6288_wire_1888);
and_n #(2, 0, 0) AND_765 (c6288_wire_1889, {c6288_wire_873_1, c6288_wire_862_1});
or_n #(2, 0, 0) OR_215 (c6288_wire_873, {c6288_wire_1814, c6288_wire_1887});
xor_n #(2, 0, 0) XOR_189 (c6288_wire_736, {c6288_wire_1890_0, c6288_wire_1891_0});
or_n #(2, 0, 0) OR_216 (c6288_wire_1890, {c6288_wire_1892, c6288_wire_1893});
and_n #(2, 0, 0) AND_766 (c6288_wire_1894, {c6288_wire_1890_1, c6288_wire_1891_1});
and_n #(2, 0, 0) AND_767 (c6288_wire_1893, {c6288_wire_1860, c6288_wire_1859_1});
notg #(0, 0) NOT_233 (c6288_wire_1892, c6288_wire_1895);
xor_n #(2, 0, 0) XOR_190 (c6288_wire_734, {c6288_wire_1896_0, c6288_wire_1897_0});
or_n #(2, 0, 0) OR_217 (c6288_wire_1896, {c6288_wire_1894, c6288_wire_1898});
and_n #(2, 0, 0) AND_768 (c6288_wire_1899, {c6288_wire_1896_1, c6288_wire_1897_1});
notg #(0, 0) NOT_234 (c6288_wire_1898, c6288_wire_1900);
xor_n #(2, 0, 0) XOR_191 (c6288_wire_732, {c6288_wire_1901_0, c6288_wire_1902_0});
or_n #(2, 0, 0) OR_218 (c6288_wire_1901, {c6288_wire_1899, c6288_wire_1903});
and_n #(2, 0, 0) AND_769 (c6288_wire_1904, {c6288_wire_1901_1, c6288_wire_1902_1});
notg #(0, 0) NOT_235 (c6288_wire_1903, c6288_wire_1905);
xor_n #(2, 0, 0) XOR_192 (c6288_wire_730, {c6288_wire_1906_0, c6288_wire_1907_0});
or_n #(2, 0, 0) OR_219 (c6288_wire_1906, {c6288_wire_1904, c6288_wire_1908});
and_n #(2, 0, 0) AND_770 (c6288_wire_1909, {c6288_wire_1906_1, c6288_wire_1907_1});
notg #(0, 0) NOT_236 (c6288_wire_1908, c6288_wire_1910);
xor_n #(2, 0, 0) XOR_193 (c6288_wire_728, {c6288_wire_1911_0, c6288_wire_1912_0});
or_n #(2, 0, 0) OR_220 (c6288_wire_1911, {c6288_wire_1909, c6288_wire_1913});
and_n #(2, 0, 0) AND_771 (c6288_wire_1914, {c6288_wire_1911_1, c6288_wire_1912_1});
notg #(0, 0) NOT_237 (c6288_wire_1913, c6288_wire_1915);
xor_n #(2, 0, 0) XOR_194 (c6288_wire_726, {c6288_wire_1916_0, c6288_wire_1917_0});
or_n #(2, 0, 0) OR_221 (c6288_wire_1916, {c6288_wire_1914, c6288_wire_1918});
and_n #(2, 0, 0) AND_772 (c6288_wire_1919, {c6288_wire_1916_1, c6288_wire_1917_1});
notg #(0, 0) NOT_238 (c6288_wire_1918, c6288_wire_1920);
xor_n #(2, 0, 0) XOR_195 (c6288_wire_724, {c6288_wire_1921_0, c6288_wire_1922_0});
or_n #(2, 0, 0) OR_222 (c6288_wire_1921, {c6288_wire_1919, c6288_wire_1923});
and_n #(2, 0, 0) AND_773 (c6288_wire_1924, {c6288_wire_1921_1, c6288_wire_1922_1});
notg #(0, 0) NOT_239 (c6288_wire_1923, c6288_wire_1925);
xor_n #(2, 0, 0) XOR_196 (c6288_wire_722, {c6288_wire_1926_0, c6288_wire_1927_0});
or_n #(2, 0, 0) OR_223 (c6288_wire_1926, {c6288_wire_1924, c6288_wire_1928});
and_n #(2, 0, 0) AND_774 (c6288_wire_1929, {c6288_wire_1926_1, c6288_wire_1927_1});
notg #(0, 0) NOT_240 (c6288_wire_1928, c6288_wire_1930);
xor_n #(2, 0, 0) XOR_197 (c6288_wire_720, {c6288_wire_1866_1, c6288_wire_1867_1});
or_n #(2, 0, 0) OR_224 (c6288_wire_1866, {c6288_wire_1929, c6288_wire_1931});
notg #(0, 0) NOT_241 (c6288_wire_1931, c6288_wire_1932);
or_n #(2, 0, 0) OR_225 (c6288_wire_1933, {c6288_wire_1934, c6288_wire_1935});
or_n #(2, 0, 0) OR_226 (c6288_wire_1936, {c6288_wire_1937, c6288_wire_1938});
or_n #(2, 0, 0) OR_227 (c6288_wire_1939, {c6288_wire_1940, c6288_wire_1941});
or_n #(2, 0, 0) OR_228 (c6288_wire_1942, {c6288_wire_1943, c6288_wire_1944});
or_n #(2, 0, 0) OR_229 (c6288_wire_1945, {c6288_wire_1946, c6288_wire_1947});
or_n #(2, 0, 0) OR_230 (c6288_wire_1948, {c6288_wire_1949, c6288_wire_1950});
or_n #(2, 0, 0) OR_231 (c6288_wire_1951, {c6288_wire_1264, c6288_wire_1952});
or_n #(2, 0, 0) OR_232 (c6288_wire_1953, {c6288_wire_1343, c6288_wire_1954});
or_n #(2, 0, 0) OR_233 (c6288_wire_1955, {c6288_wire_1956, c6288_wire_34});
or_n #(2, 0, 0) OR_234 (c6288_wire_1957, {c6288_wire_1421, c6288_wire_1958});
or_n #(2, 0, 0) OR_235 (c6288_wire_1959, {c6288_wire_1499, c6288_wire_1960});
or_n #(2, 0, 0) OR_236 (c6288_wire_1961, {c6288_wire_1577, c6288_wire_1962});
or_n #(2, 0, 0) OR_237 (c6288_wire_1963, {c6288_wire_1655, c6288_wire_1964});
or_n #(2, 0, 0) OR_238 (c6288_wire_1965, {c6288_wire_1733, c6288_wire_1966});
or_n #(2, 0, 0) OR_239 (c6288_wire_1967, {c6288_wire_1811, c6288_wire_1968});
or_n #(2, 0, 0) OR_240 (c6288_wire_1969, {c6288_wire_1889, c6288_wire_1970});
or_n #(2, 0, 0) OR_241 (c6288_wire_1971, {c6288_wire_868, c6288_wire_1972});
or_n #(2, 0, 0) OR_242 (c6288_wire_1973, {c6288_wire_948, c6288_wire_1974});
or_n #(2, 0, 0) OR_243 (c6288_wire_1975, {c6288_wire_1026, c6288_wire_1976});
or_n #(2, 0, 0) OR_244 (c6288_wire_1977, {c6288_wire_1978, c6288_wire_1979});
or_n #(2, 0, 0) OR_245 (c6288_wire_1980, {c6288_wire_1102, c6288_wire_1981});
or_n #(2, 0, 0) OR_246 (c6288_wire_1982, {c6288_wire_1983, c6288_wire_1984});
or_n #(2, 0, 0) OR_247 (c6288_wire_1985, {c6288_wire_1986, c6288_wire_1987});
or_n #(2, 0, 0) OR_248 (c6288_wire_1988, {c6288_wire_1989, c6288_wire_1990});
or_n #(2, 0, 0) OR_249 (c6288_wire_1991, {c6288_wire_1992, c6288_wire_1993});
or_n #(2, 0, 0) OR_250 (c6288_wire_1994, {c6288_wire_1995, c6288_wire_1996});
or_n #(2, 0, 0) OR_251 (c6288_wire_1997, {c6288_wire_1998, c6288_wire_1999});
or_n #(2, 0, 0) OR_252 (c6288_wire_2000, {c6288_wire_2001, c6288_wire_2002});
nand_n #(2, 0, 0) NAND_1 (c6288_wire_35, {c6288_wire_32_31, c6288_wire_6_32});
and_n #(2, 0, 0) AND_775 (c6288_wire_1956, {c6288_wire_76, c6288_wire_33});
notg #(0, 0) NOT_242 (c6288_wire_2003, c6288_wire_756_1);
and_n #(2, 0, 0) AND_776 (c6288_wire_1937, {c6288_wire_2003, c6288_wire_833_0});
and_n #(2, 0, 0) AND_777 (c6288_wire_1938, {c6288_wire_106, c6288_wire_2004});
notg #(0, 0) NOT_243 (c6288_wire_2004, c6288_wire_833_1);
and_n #(2, 0, 0) AND_778 (c6288_wire_1978, {c6288_wire_79, c6288_wire_2005});
notg #(0, 0) NOT_244 (c6288_wire_2006, c6288_wire_762_1);
and_n #(2, 0, 0) AND_779 (c6288_wire_1940, {c6288_wire_2006, c6288_wire_748_0});
and_n #(2, 0, 0) AND_780 (c6288_wire_1941, {c6288_wire_109, c6288_wire_2007});
notg #(0, 0) NOT_245 (c6288_wire_2007, c6288_wire_748_1);
notg #(0, 0) NOT_246 (c6288_wire_2008, c6288_wire_768_1);
and_n #(2, 0, 0) AND_781 (c6288_wire_1943, {c6288_wire_2008, c6288_wire_757_0});
and_n #(2, 0, 0) AND_782 (c6288_wire_1944, {c6288_wire_112, c6288_wire_2009});
notg #(0, 0) NOT_247 (c6288_wire_2009, c6288_wire_757_1);
notg #(0, 0) NOT_248 (c6288_wire_2010, c6288_wire_774_1);
and_n #(2, 0, 0) AND_783 (c6288_wire_1946, {c6288_wire_2010, c6288_wire_763_0});
and_n #(2, 0, 0) AND_784 (c6288_wire_1947, {c6288_wire_115, c6288_wire_2011});
notg #(0, 0) NOT_249 (c6288_wire_2011, c6288_wire_763_1);
notg #(0, 0) NOT_250 (c6288_wire_2012, c6288_wire_779_1);
and_n #(2, 0, 0) AND_785 (c6288_wire_1949, {c6288_wire_2012, c6288_wire_769_0});
and_n #(2, 0, 0) AND_786 (c6288_wire_1950, {c6288_wire_118, c6288_wire_2013});
notg #(0, 0) NOT_251 (c6288_wire_2013, c6288_wire_769_1);
notg #(0, 0) NOT_252 (c6288_wire_2014, c6288_wire_790_1);
and_n #(2, 0, 0) AND_787 (c6288_wire_1979, {c6288_wire_2014, c6288_wire_2015_0});
notg #(0, 0) NOT_253 (c6288_wire_2005, c6288_wire_2015_1);
notg #(0, 0) NOT_254 (c6288_wire_2016, c6288_wire_796_1);
and_n #(2, 0, 0) AND_788 (c6288_wire_1983, {c6288_wire_2016, c6288_wire_784_0});
and_n #(2, 0, 0) AND_789 (c6288_wire_1984, {c6288_wire_82, c6288_wire_2017});
notg #(0, 0) NOT_255 (c6288_wire_2017, c6288_wire_784_1);
notg #(0, 0) NOT_256 (c6288_wire_2018, c6288_wire_802_1);
and_n #(2, 0, 0) AND_790 (c6288_wire_1986, {c6288_wire_2018, c6288_wire_791_0});
and_n #(2, 0, 0) AND_791 (c6288_wire_1987, {c6288_wire_85, c6288_wire_2019});
notg #(0, 0) NOT_257 (c6288_wire_2019, c6288_wire_791_1);
notg #(0, 0) NOT_258 (c6288_wire_2020, c6288_wire_808_1);
and_n #(2, 0, 0) AND_792 (c6288_wire_1989, {c6288_wire_2020, c6288_wire_797_0});
and_n #(2, 0, 0) AND_793 (c6288_wire_1990, {c6288_wire_88, c6288_wire_2021});
notg #(0, 0) NOT_259 (c6288_wire_2021, c6288_wire_797_1);
notg #(0, 0) NOT_260 (c6288_wire_2022, c6288_wire_814_1);
and_n #(2, 0, 0) AND_794 (c6288_wire_1992, {c6288_wire_2022, c6288_wire_803_0});
and_n #(2, 0, 0) AND_795 (c6288_wire_1993, {c6288_wire_91, c6288_wire_2023});
notg #(0, 0) NOT_261 (c6288_wire_2023, c6288_wire_803_1);
notg #(0, 0) NOT_262 (c6288_wire_2024, c6288_wire_820_1);
and_n #(2, 0, 0) AND_796 (c6288_wire_1995, {c6288_wire_2024, c6288_wire_809_0});
and_n #(2, 0, 0) AND_797 (c6288_wire_1996, {c6288_wire_94, c6288_wire_2025});
notg #(0, 0) NOT_263 (c6288_wire_2025, c6288_wire_809_1);
notg #(0, 0) NOT_264 (c6288_wire_2026, c6288_wire_826_1);
and_n #(2, 0, 0) AND_798 (c6288_wire_1998, {c6288_wire_2026, c6288_wire_815_0});
and_n #(2, 0, 0) AND_799 (c6288_wire_1999, {c6288_wire_97, c6288_wire_2027});
notg #(0, 0) NOT_265 (c6288_wire_2027, c6288_wire_815_1);
notg #(0, 0) NOT_266 (c6288_wire_2028, c6288_wire_832_1);
and_n #(2, 0, 0) AND_800 (c6288_wire_2001, {c6288_wire_2028, c6288_wire_821_0});
and_n #(2, 0, 0) AND_801 (c6288_wire_2002, {c6288_wire_100, c6288_wire_2029});
notg #(0, 0) NOT_267 (c6288_wire_2029, c6288_wire_821_1);
notg #(0, 0) NOT_268 (c6288_wire_2030, c6288_wire_835_1);
and_n #(2, 0, 0) AND_802 (c6288_wire_1934, {c6288_wire_2030, c6288_wire_827_0});
and_n #(2, 0, 0) AND_803 (c6288_wire_1935, {c6288_wire_103, c6288_wire_2031});
notg #(0, 0) NOT_269 (c6288_wire_2031, c6288_wire_827_1);
or_n #(2, 0, 0) OR_253 (c6288_wire_1859, {c6288_wire_13, c6288_wire_2032});
nand_n #(2, 0, 0) NAND_2 (c6288_wire_2033, {c6288_wire_2_31, c6288_wire_6_33});
and_n #(2, 0, 0) AND_804 (c6288_wire_2032, {c6288_wire_12, c6288_wire_2033});
or_n #(2, 0, 0) OR_254 (c6288_wire_1862, {c6288_wire_141, c6288_wire_2034});
nand_n #(2, 0, 0) NAND_3 (c6288_wire_2035, {c6288_wire_2_32, c6288_wire_105_32});
notg #(0, 0) NOT_270 (c6288_wire_2036, c6288_wire_142_1);
and_n #(2, 0, 0) AND_805 (c6288_wire_2034, {c6288_wire_2036, c6288_wire_2035});
or_n #(2, 0, 0) OR_255 (c6288_wire_1870, {c6288_wire_139, c6288_wire_2037});
nand_n #(2, 0, 0) NAND_4 (c6288_wire_2038, {c6288_wire_2_33, c6288_wire_108_32});
notg #(0, 0) NOT_271 (c6288_wire_2039, c6288_wire_140_1);
and_n #(2, 0, 0) AND_806 (c6288_wire_2037, {c6288_wire_2039, c6288_wire_2038});
or_n #(2, 0, 0) OR_256 (c6288_wire_1875, {c6288_wire_137, c6288_wire_2040});
nand_n #(2, 0, 0) NAND_5 (c6288_wire_2041, {c6288_wire_2_34, c6288_wire_111_32});
notg #(0, 0) NOT_272 (c6288_wire_2042, c6288_wire_138_1);
and_n #(2, 0, 0) AND_807 (c6288_wire_2040, {c6288_wire_2042, c6288_wire_2041});
or_n #(2, 0, 0) OR_257 (c6288_wire_1880, {c6288_wire_135, c6288_wire_2043});
nand_n #(2, 0, 0) NAND_6 (c6288_wire_2044, {c6288_wire_2_35, c6288_wire_114_32});
notg #(0, 0) NOT_273 (c6288_wire_2045, c6288_wire_136_1);
and_n #(2, 0, 0) AND_808 (c6288_wire_2043, {c6288_wire_2045, c6288_wire_2044});
or_n #(2, 0, 0) OR_258 (c6288_wire_1885, {c6288_wire_133, c6288_wire_2046});
nand_n #(2, 0, 0) NAND_7 (c6288_wire_2047, {c6288_wire_2_36, c6288_wire_117_32});
notg #(0, 0) NOT_274 (c6288_wire_2048, c6288_wire_134_1);
and_n #(2, 0, 0) AND_809 (c6288_wire_2046, {c6288_wire_2048, c6288_wire_2047});
nor_n #(2, 0, 0) NOR_3 (c6288_wire_1970, {c6288_wire_862_2, c6288_wire_873_2});
or_n #(2, 0, 0) OR_259 (c6288_wire_1891, {c6288_wire_159, c6288_wire_2049});
nand_n #(2, 0, 0) NAND_8 (c6288_wire_2050, {c6288_wire_2_37, c6288_wire_78_33});
notg #(0, 0) NOT_275 (c6288_wire_2051, c6288_wire_160_1);
and_n #(2, 0, 0) AND_810 (c6288_wire_2049, {c6288_wire_2051, c6288_wire_2050});
or_n #(2, 0, 0) OR_260 (c6288_wire_1897, {c6288_wire_157, c6288_wire_2052});
nand_n #(2, 0, 0) NAND_9 (c6288_wire_2053, {c6288_wire_2_38, c6288_wire_81_32});
notg #(0, 0) NOT_276 (c6288_wire_2054, c6288_wire_158_1);
and_n #(2, 0, 0) AND_811 (c6288_wire_2052, {c6288_wire_2054, c6288_wire_2053});
or_n #(2, 0, 0) OR_261 (c6288_wire_1902, {c6288_wire_155, c6288_wire_2055});
nand_n #(2, 0, 0) NAND_10 (c6288_wire_2056, {c6288_wire_2_39, c6288_wire_84_32});
notg #(0, 0) NOT_277 (c6288_wire_2057, c6288_wire_156_1);
and_n #(2, 0, 0) AND_812 (c6288_wire_2055, {c6288_wire_2057, c6288_wire_2056});
or_n #(2, 0, 0) OR_262 (c6288_wire_1907, {c6288_wire_153, c6288_wire_2058});
nand_n #(2, 0, 0) NAND_11 (c6288_wire_2059, {c6288_wire_2_40, c6288_wire_87_32});
notg #(0, 0) NOT_278 (c6288_wire_2060, c6288_wire_154_1);
and_n #(2, 0, 0) AND_813 (c6288_wire_2058, {c6288_wire_2060, c6288_wire_2059});
or_n #(2, 0, 0) OR_263 (c6288_wire_1912, {c6288_wire_151, c6288_wire_2061});
nand_n #(2, 0, 0) NAND_12 (c6288_wire_2062, {c6288_wire_2_41, c6288_wire_90_32});
notg #(0, 0) NOT_279 (c6288_wire_2063, c6288_wire_152_1);
and_n #(2, 0, 0) AND_814 (c6288_wire_2061, {c6288_wire_2063, c6288_wire_2062});
or_n #(2, 0, 0) OR_264 (c6288_wire_1917, {c6288_wire_149, c6288_wire_2064});
nand_n #(2, 0, 0) NAND_13 (c6288_wire_2065, {c6288_wire_2_42, c6288_wire_93_32});
notg #(0, 0) NOT_280 (c6288_wire_2066, c6288_wire_150_1);
and_n #(2, 0, 0) AND_815 (c6288_wire_2064, {c6288_wire_2066, c6288_wire_2065});
or_n #(2, 0, 0) OR_265 (c6288_wire_1922, {c6288_wire_147, c6288_wire_2067});
nand_n #(2, 0, 0) NAND_14 (c6288_wire_2068, {c6288_wire_2_43, c6288_wire_96_32});
notg #(0, 0) NOT_281 (c6288_wire_2069, c6288_wire_148_1);
and_n #(2, 0, 0) AND_816 (c6288_wire_2067, {c6288_wire_2069, c6288_wire_2068});
or_n #(2, 0, 0) OR_266 (c6288_wire_1927, {c6288_wire_145, c6288_wire_2070});
nand_n #(2, 0, 0) NAND_15 (c6288_wire_2071, {c6288_wire_2_44, c6288_wire_99_32});
notg #(0, 0) NOT_282 (c6288_wire_2072, c6288_wire_146_1);
and_n #(2, 0, 0) AND_817 (c6288_wire_2070, {c6288_wire_2072, c6288_wire_2071});
or_n #(2, 0, 0) OR_267 (c6288_wire_1867, {c6288_wire_143, c6288_wire_2073});
nand_n #(2, 0, 0) NAND_16 (c6288_wire_2074, {c6288_wire_2_45, c6288_wire_102_32});
notg #(0, 0) NOT_283 (c6288_wire_2075, c6288_wire_144_1);
and_n #(2, 0, 0) AND_818 (c6288_wire_2073, {c6288_wire_2075, c6288_wire_2074});
or_n #(2, 0, 0) OR_268 (c6288_wire_837, {c6288_wire_18, c6288_wire_2076});
nand_n #(2, 0, 0) NAND_17 (c6288_wire_2077, {c6288_wire_10_31, c6288_wire_6_34});
and_n #(2, 0, 0) AND_819 (c6288_wire_2076, {c6288_wire_17, c6288_wire_2077});
or_n #(2, 0, 0) OR_269 (c6288_wire_840, {c6288_wire_183, c6288_wire_2078});
nand_n #(2, 0, 0) NAND_18 (c6288_wire_2079, {c6288_wire_10_32, c6288_wire_105_33});
notg #(0, 0) NOT_284 (c6288_wire_2080, c6288_wire_184_1);
and_n #(2, 0, 0) AND_820 (c6288_wire_2078, {c6288_wire_2080, c6288_wire_2079});
or_n #(2, 0, 0) OR_270 (c6288_wire_848, {c6288_wire_181, c6288_wire_2081});
nand_n #(2, 0, 0) NAND_19 (c6288_wire_2082, {c6288_wire_10_33, c6288_wire_108_33});
notg #(0, 0) NOT_285 (c6288_wire_2083, c6288_wire_182_1);
and_n #(2, 0, 0) AND_821 (c6288_wire_2081, {c6288_wire_2083, c6288_wire_2082});
or_n #(2, 0, 0) OR_271 (c6288_wire_853, {c6288_wire_179, c6288_wire_2084});
nand_n #(2, 0, 0) NAND_20 (c6288_wire_2085, {c6288_wire_10_34, c6288_wire_111_33});
notg #(0, 0) NOT_286 (c6288_wire_2086, c6288_wire_180_1);
and_n #(2, 0, 0) AND_822 (c6288_wire_2084, {c6288_wire_2086, c6288_wire_2085});
or_n #(2, 0, 0) OR_272 (c6288_wire_858, {c6288_wire_177, c6288_wire_2087});
nand_n #(2, 0, 0) NAND_21 (c6288_wire_2088, {c6288_wire_10_35, c6288_wire_114_33});
notg #(0, 0) NOT_287 (c6288_wire_2089, c6288_wire_178_1);
and_n #(2, 0, 0) AND_823 (c6288_wire_2087, {c6288_wire_2089, c6288_wire_2088});
or_n #(2, 0, 0) OR_273 (c6288_wire_864, {c6288_wire_175, c6288_wire_2090});
nand_n #(2, 0, 0) NAND_22 (c6288_wire_2091, {c6288_wire_10_36, c6288_wire_117_33});
notg #(0, 0) NOT_288 (c6288_wire_2092, c6288_wire_176_1);
and_n #(2, 0, 0) AND_824 (c6288_wire_2090, {c6288_wire_2092, c6288_wire_2091});
nor_n #(2, 0, 0) NOR_4 (c6288_wire_1972, {c6288_wire_870_2, c6288_wire_869_2});
or_n #(2, 0, 0) OR_274 (c6288_wire_875, {c6288_wire_201, c6288_wire_2093});
nand_n #(2, 0, 0) NAND_23 (c6288_wire_2094, {c6288_wire_10_37, c6288_wire_78_34});
notg #(0, 0) NOT_289 (c6288_wire_2095, c6288_wire_202_1);
and_n #(2, 0, 0) AND_825 (c6288_wire_2093, {c6288_wire_2095, c6288_wire_2094});
or_n #(2, 0, 0) OR_275 (c6288_wire_881, {c6288_wire_199, c6288_wire_2096});
nand_n #(2, 0, 0) NAND_24 (c6288_wire_2097, {c6288_wire_10_38, c6288_wire_81_33});
notg #(0, 0) NOT_290 (c6288_wire_2098, c6288_wire_200_1);
and_n #(2, 0, 0) AND_826 (c6288_wire_2096, {c6288_wire_2098, c6288_wire_2097});
or_n #(2, 0, 0) OR_276 (c6288_wire_886, {c6288_wire_197, c6288_wire_2099});
nand_n #(2, 0, 0) NAND_25 (c6288_wire_2100, {c6288_wire_10_39, c6288_wire_84_33});
notg #(0, 0) NOT_291 (c6288_wire_2101, c6288_wire_198_1);
and_n #(2, 0, 0) AND_827 (c6288_wire_2099, {c6288_wire_2101, c6288_wire_2100});
or_n #(2, 0, 0) OR_277 (c6288_wire_891, {c6288_wire_195, c6288_wire_2102});
nand_n #(2, 0, 0) NAND_26 (c6288_wire_2103, {c6288_wire_10_40, c6288_wire_87_33});
notg #(0, 0) NOT_292 (c6288_wire_2104, c6288_wire_196_1);
and_n #(2, 0, 0) AND_828 (c6288_wire_2102, {c6288_wire_2104, c6288_wire_2103});
or_n #(2, 0, 0) OR_278 (c6288_wire_896, {c6288_wire_193, c6288_wire_2105});
nand_n #(2, 0, 0) NAND_27 (c6288_wire_2106, {c6288_wire_10_41, c6288_wire_90_33});
notg #(0, 0) NOT_293 (c6288_wire_2107, c6288_wire_194_1);
and_n #(2, 0, 0) AND_829 (c6288_wire_2105, {c6288_wire_2107, c6288_wire_2106});
or_n #(2, 0, 0) OR_279 (c6288_wire_901, {c6288_wire_191, c6288_wire_2108});
nand_n #(2, 0, 0) NAND_28 (c6288_wire_2109, {c6288_wire_10_42, c6288_wire_93_33});
notg #(0, 0) NOT_294 (c6288_wire_2110, c6288_wire_192_1);
and_n #(2, 0, 0) AND_830 (c6288_wire_2108, {c6288_wire_2110, c6288_wire_2109});
or_n #(2, 0, 0) OR_280 (c6288_wire_906, {c6288_wire_189, c6288_wire_2111});
nand_n #(2, 0, 0) NAND_29 (c6288_wire_2112, {c6288_wire_10_43, c6288_wire_96_33});
notg #(0, 0) NOT_295 (c6288_wire_2113, c6288_wire_190_1);
and_n #(2, 0, 0) AND_831 (c6288_wire_2111, {c6288_wire_2113, c6288_wire_2112});
or_n #(2, 0, 0) OR_281 (c6288_wire_911, {c6288_wire_187, c6288_wire_2114});
nand_n #(2, 0, 0) NAND_30 (c6288_wire_2115, {c6288_wire_10_44, c6288_wire_99_33});
notg #(0, 0) NOT_296 (c6288_wire_2116, c6288_wire_188_1);
and_n #(2, 0, 0) AND_832 (c6288_wire_2114, {c6288_wire_2116, c6288_wire_2115});
or_n #(2, 0, 0) OR_282 (c6288_wire_845, {c6288_wire_185, c6288_wire_2117});
nand_n #(2, 0, 0) NAND_31 (c6288_wire_2118, {c6288_wire_10_45, c6288_wire_102_33});
notg #(0, 0) NOT_297 (c6288_wire_2119, c6288_wire_186_1);
and_n #(2, 0, 0) AND_833 (c6288_wire_2117, {c6288_wire_2119, c6288_wire_2118});
or_n #(2, 0, 0) OR_283 (c6288_wire_918, {c6288_wire_23, c6288_wire_2120});
nand_n #(2, 0, 0) NAND_32 (c6288_wire_2121, {c6288_wire_15_31, c6288_wire_6_35});
and_n #(2, 0, 0) AND_834 (c6288_wire_2120, {c6288_wire_22, c6288_wire_2121});
or_n #(2, 0, 0) OR_284 (c6288_wire_921, {c6288_wire_225, c6288_wire_2122});
nand_n #(2, 0, 0) NAND_33 (c6288_wire_2123, {c6288_wire_15_32, c6288_wire_105_34});
notg #(0, 0) NOT_298 (c6288_wire_2124, c6288_wire_226_1);
and_n #(2, 0, 0) AND_835 (c6288_wire_2122, {c6288_wire_2124, c6288_wire_2123});
or_n #(2, 0, 0) OR_285 (c6288_wire_929, {c6288_wire_223, c6288_wire_2125});
nand_n #(2, 0, 0) NAND_34 (c6288_wire_2126, {c6288_wire_15_33, c6288_wire_108_34});
notg #(0, 0) NOT_299 (c6288_wire_2127, c6288_wire_224_1);
and_n #(2, 0, 0) AND_836 (c6288_wire_2125, {c6288_wire_2127, c6288_wire_2126});
or_n #(2, 0, 0) OR_286 (c6288_wire_934, {c6288_wire_221, c6288_wire_2128});
nand_n #(2, 0, 0) NAND_35 (c6288_wire_2129, {c6288_wire_15_34, c6288_wire_111_34});
notg #(0, 0) NOT_300 (c6288_wire_2130, c6288_wire_222_1);
and_n #(2, 0, 0) AND_837 (c6288_wire_2128, {c6288_wire_2130, c6288_wire_2129});
or_n #(2, 0, 0) OR_287 (c6288_wire_939, {c6288_wire_219, c6288_wire_2131});
nand_n #(2, 0, 0) NAND_36 (c6288_wire_2132, {c6288_wire_15_35, c6288_wire_114_34});
notg #(0, 0) NOT_301 (c6288_wire_2133, c6288_wire_220_1);
and_n #(2, 0, 0) AND_838 (c6288_wire_2131, {c6288_wire_2133, c6288_wire_2132});
or_n #(2, 0, 0) OR_288 (c6288_wire_944, {c6288_wire_217, c6288_wire_2134});
nand_n #(2, 0, 0) NAND_37 (c6288_wire_2135, {c6288_wire_15_36, c6288_wire_117_34});
notg #(0, 0) NOT_302 (c6288_wire_2136, c6288_wire_218_1);
and_n #(2, 0, 0) AND_839 (c6288_wire_2134, {c6288_wire_2136, c6288_wire_2135});
nor_n #(2, 0, 0) NOR_5 (c6288_wire_1974, {c6288_wire_950_2, c6288_wire_949_2});
or_n #(2, 0, 0) OR_289 (c6288_wire_953, {c6288_wire_243, c6288_wire_2137});
nand_n #(2, 0, 0) NAND_38 (c6288_wire_2138, {c6288_wire_15_37, c6288_wire_78_35});
notg #(0, 0) NOT_303 (c6288_wire_2139, c6288_wire_244_1);
and_n #(2, 0, 0) AND_840 (c6288_wire_2137, {c6288_wire_2139, c6288_wire_2138});
or_n #(2, 0, 0) OR_290 (c6288_wire_959, {c6288_wire_241, c6288_wire_2140});
nand_n #(2, 0, 0) NAND_39 (c6288_wire_2141, {c6288_wire_15_38, c6288_wire_81_34});
notg #(0, 0) NOT_304 (c6288_wire_2142, c6288_wire_242_1);
and_n #(2, 0, 0) AND_841 (c6288_wire_2140, {c6288_wire_2142, c6288_wire_2141});
or_n #(2, 0, 0) OR_291 (c6288_wire_964, {c6288_wire_239, c6288_wire_2143});
nand_n #(2, 0, 0) NAND_40 (c6288_wire_2144, {c6288_wire_15_39, c6288_wire_84_34});
notg #(0, 0) NOT_305 (c6288_wire_2145, c6288_wire_240_1);
and_n #(2, 0, 0) AND_842 (c6288_wire_2143, {c6288_wire_2145, c6288_wire_2144});
or_n #(2, 0, 0) OR_292 (c6288_wire_969, {c6288_wire_237, c6288_wire_2146});
nand_n #(2, 0, 0) NAND_41 (c6288_wire_2147, {c6288_wire_15_40, c6288_wire_87_34});
notg #(0, 0) NOT_306 (c6288_wire_2148, c6288_wire_238_1);
and_n #(2, 0, 0) AND_843 (c6288_wire_2146, {c6288_wire_2148, c6288_wire_2147});
or_n #(2, 0, 0) OR_293 (c6288_wire_974, {c6288_wire_235, c6288_wire_2149});
nand_n #(2, 0, 0) NAND_42 (c6288_wire_2150, {c6288_wire_15_41, c6288_wire_90_34});
notg #(0, 0) NOT_307 (c6288_wire_2151, c6288_wire_236_1);
and_n #(2, 0, 0) AND_844 (c6288_wire_2149, {c6288_wire_2151, c6288_wire_2150});
or_n #(2, 0, 0) OR_294 (c6288_wire_979, {c6288_wire_233, c6288_wire_2152});
nand_n #(2, 0, 0) NAND_43 (c6288_wire_2153, {c6288_wire_15_42, c6288_wire_93_34});
notg #(0, 0) NOT_308 (c6288_wire_2154, c6288_wire_234_1);
and_n #(2, 0, 0) AND_845 (c6288_wire_2152, {c6288_wire_2154, c6288_wire_2153});
or_n #(2, 0, 0) OR_295 (c6288_wire_984, {c6288_wire_231, c6288_wire_2155});
nand_n #(2, 0, 0) NAND_44 (c6288_wire_2156, {c6288_wire_15_43, c6288_wire_96_34});
notg #(0, 0) NOT_309 (c6288_wire_2157, c6288_wire_232_1);
and_n #(2, 0, 0) AND_846 (c6288_wire_2155, {c6288_wire_2157, c6288_wire_2156});
or_n #(2, 0, 0) OR_296 (c6288_wire_989, {c6288_wire_229, c6288_wire_2158});
nand_n #(2, 0, 0) NAND_45 (c6288_wire_2159, {c6288_wire_15_44, c6288_wire_99_34});
notg #(0, 0) NOT_310 (c6288_wire_2160, c6288_wire_230_1);
and_n #(2, 0, 0) AND_847 (c6288_wire_2158, {c6288_wire_2160, c6288_wire_2159});
or_n #(2, 0, 0) OR_297 (c6288_wire_926, {c6288_wire_227, c6288_wire_2161});
nand_n #(2, 0, 0) NAND_46 (c6288_wire_2162, {c6288_wire_15_45, c6288_wire_102_34});
notg #(0, 0) NOT_311 (c6288_wire_2163, c6288_wire_228_1);
and_n #(2, 0, 0) AND_848 (c6288_wire_2161, {c6288_wire_2163, c6288_wire_2162});
or_n #(2, 0, 0) OR_298 (c6288_wire_996, {c6288_wire_28, c6288_wire_2164});
nand_n #(2, 0, 0) NAND_47 (c6288_wire_2165, {c6288_wire_20_31, c6288_wire_6_36});
and_n #(2, 0, 0) AND_849 (c6288_wire_2164, {c6288_wire_27, c6288_wire_2165});
or_n #(2, 0, 0) OR_299 (c6288_wire_999, {c6288_wire_267, c6288_wire_2166});
nand_n #(2, 0, 0) NAND_48 (c6288_wire_2167, {c6288_wire_20_32, c6288_wire_105_35});
notg #(0, 0) NOT_312 (c6288_wire_2168, c6288_wire_268_1);
and_n #(2, 0, 0) AND_850 (c6288_wire_2166, {c6288_wire_2168, c6288_wire_2167});
or_n #(2, 0, 0) OR_300 (c6288_wire_1007, {c6288_wire_265, c6288_wire_2169});
nand_n #(2, 0, 0) NAND_49 (c6288_wire_2170, {c6288_wire_20_33, c6288_wire_108_35});
notg #(0, 0) NOT_313 (c6288_wire_2171, c6288_wire_266_1);
and_n #(2, 0, 0) AND_851 (c6288_wire_2169, {c6288_wire_2171, c6288_wire_2170});
or_n #(2, 0, 0) OR_301 (c6288_wire_1012, {c6288_wire_263, c6288_wire_2172});
nand_n #(2, 0, 0) NAND_50 (c6288_wire_2173, {c6288_wire_20_34, c6288_wire_111_35});
notg #(0, 0) NOT_314 (c6288_wire_2174, c6288_wire_264_1);
and_n #(2, 0, 0) AND_852 (c6288_wire_2172, {c6288_wire_2174, c6288_wire_2173});
or_n #(2, 0, 0) OR_302 (c6288_wire_1017, {c6288_wire_261, c6288_wire_2175});
nand_n #(2, 0, 0) NAND_51 (c6288_wire_2176, {c6288_wire_20_35, c6288_wire_114_35});
notg #(0, 0) NOT_315 (c6288_wire_2177, c6288_wire_262_1);
and_n #(2, 0, 0) AND_853 (c6288_wire_2175, {c6288_wire_2177, c6288_wire_2176});
or_n #(2, 0, 0) OR_303 (c6288_wire_1022, {c6288_wire_259, c6288_wire_2178});
nand_n #(2, 0, 0) NAND_52 (c6288_wire_2179, {c6288_wire_20_36, c6288_wire_117_35});
notg #(0, 0) NOT_316 (c6288_wire_2180, c6288_wire_260_1);
and_n #(2, 0, 0) AND_854 (c6288_wire_2178, {c6288_wire_2180, c6288_wire_2179});
nor_n #(2, 0, 0) NOR_6 (c6288_wire_1976, {c6288_wire_1028_2, c6288_wire_1027_2});
or_n #(2, 0, 0) OR_304 (c6288_wire_1031, {c6288_wire_285, c6288_wire_2181});
nand_n #(2, 0, 0) NAND_53 (c6288_wire_2182, {c6288_wire_20_37, c6288_wire_78_36});
notg #(0, 0) NOT_317 (c6288_wire_2183, c6288_wire_286_1);
and_n #(2, 0, 0) AND_855 (c6288_wire_2181, {c6288_wire_2183, c6288_wire_2182});
or_n #(2, 0, 0) OR_305 (c6288_wire_1037, {c6288_wire_283, c6288_wire_2184});
nand_n #(2, 0, 0) NAND_54 (c6288_wire_2185, {c6288_wire_20_38, c6288_wire_81_35});
notg #(0, 0) NOT_318 (c6288_wire_2186, c6288_wire_284_1);
and_n #(2, 0, 0) AND_856 (c6288_wire_2184, {c6288_wire_2186, c6288_wire_2185});
or_n #(2, 0, 0) OR_306 (c6288_wire_1042, {c6288_wire_281, c6288_wire_2187});
nand_n #(2, 0, 0) NAND_55 (c6288_wire_2188, {c6288_wire_20_39, c6288_wire_84_35});
notg #(0, 0) NOT_319 (c6288_wire_2189, c6288_wire_282_1);
and_n #(2, 0, 0) AND_857 (c6288_wire_2187, {c6288_wire_2189, c6288_wire_2188});
or_n #(2, 0, 0) OR_307 (c6288_wire_1047, {c6288_wire_279, c6288_wire_2190});
nand_n #(2, 0, 0) NAND_56 (c6288_wire_2191, {c6288_wire_20_40, c6288_wire_87_35});
notg #(0, 0) NOT_320 (c6288_wire_2192, c6288_wire_280_1);
and_n #(2, 0, 0) AND_858 (c6288_wire_2190, {c6288_wire_2192, c6288_wire_2191});
or_n #(2, 0, 0) OR_308 (c6288_wire_1052, {c6288_wire_277, c6288_wire_2193});
nand_n #(2, 0, 0) NAND_57 (c6288_wire_2194, {c6288_wire_20_41, c6288_wire_90_35});
notg #(0, 0) NOT_321 (c6288_wire_2195, c6288_wire_278_1);
and_n #(2, 0, 0) AND_859 (c6288_wire_2193, {c6288_wire_2195, c6288_wire_2194});
or_n #(2, 0, 0) OR_309 (c6288_wire_1057, {c6288_wire_275, c6288_wire_2196});
nand_n #(2, 0, 0) NAND_58 (c6288_wire_2197, {c6288_wire_20_42, c6288_wire_93_35});
notg #(0, 0) NOT_322 (c6288_wire_2198, c6288_wire_276_1);
and_n #(2, 0, 0) AND_860 (c6288_wire_2196, {c6288_wire_2198, c6288_wire_2197});
or_n #(2, 0, 0) OR_310 (c6288_wire_1062, {c6288_wire_273, c6288_wire_2199});
nand_n #(2, 0, 0) NAND_59 (c6288_wire_2200, {c6288_wire_20_43, c6288_wire_96_35});
notg #(0, 0) NOT_323 (c6288_wire_2201, c6288_wire_274_1);
and_n #(2, 0, 0) AND_861 (c6288_wire_2199, {c6288_wire_2201, c6288_wire_2200});
or_n #(2, 0, 0) OR_311 (c6288_wire_1067, {c6288_wire_271, c6288_wire_2202});
nand_n #(2, 0, 0) NAND_60 (c6288_wire_2203, {c6288_wire_20_44, c6288_wire_99_35});
notg #(0, 0) NOT_324 (c6288_wire_2204, c6288_wire_272_1);
and_n #(2, 0, 0) AND_862 (c6288_wire_2202, {c6288_wire_2204, c6288_wire_2203});
or_n #(2, 0, 0) OR_312 (c6288_wire_1004, {c6288_wire_269, c6288_wire_2205});
nand_n #(2, 0, 0) NAND_61 (c6288_wire_2206, {c6288_wire_20_45, c6288_wire_102_35});
notg #(0, 0) NOT_325 (c6288_wire_2207, c6288_wire_270_1);
and_n #(2, 0, 0) AND_863 (c6288_wire_2205, {c6288_wire_2207, c6288_wire_2206});
or_n #(2, 0, 0) OR_313 (c6288_wire_1073, {c6288_wire_2208, c6288_wire_2209});
and_n #(2, 0, 0) AND_864 (c6288_wire_2209, {c6288_wire_328, c6288_wire_2210});
and_n #(2, 0, 0) AND_865 (c6288_wire_2208, {c6288_wire_356, c6288_wire_2211});
nand_n #(2, 0, 0) NAND_62 (c6288_wire_2210, {c6288_wire_330_30, c6288_wire_3_16});
nand_n #(2, 0, 0) NAND_63 (c6288_wire_2211, {c6288_wire_25_30, c6288_wire_6_37});
or_n #(2, 0, 0) OR_314 (c6288_wire_1075, {c6288_wire_310, c6288_wire_2212});
nand_n #(2, 0, 0) NAND_64 (c6288_wire_2213, {c6288_wire_25_31, c6288_wire_105_36});
notg #(0, 0) NOT_326 (c6288_wire_2214, c6288_wire_311_1);
and_n #(2, 0, 0) AND_866 (c6288_wire_2212, {c6288_wire_2214, c6288_wire_2213});
or_n #(2, 0, 0) OR_315 (c6288_wire_1083, {c6288_wire_308, c6288_wire_2215});
nand_n #(2, 0, 0) NAND_65 (c6288_wire_2216, {c6288_wire_25_32, c6288_wire_108_36});
notg #(0, 0) NOT_327 (c6288_wire_2217, c6288_wire_309_1);
and_n #(2, 0, 0) AND_867 (c6288_wire_2215, {c6288_wire_2217, c6288_wire_2216});
or_n #(2, 0, 0) OR_316 (c6288_wire_1088, {c6288_wire_306, c6288_wire_2218});
nand_n #(2, 0, 0) NAND_66 (c6288_wire_2219, {c6288_wire_25_33, c6288_wire_111_36});
notg #(0, 0) NOT_328 (c6288_wire_2220, c6288_wire_307_1);
and_n #(2, 0, 0) AND_868 (c6288_wire_2218, {c6288_wire_2220, c6288_wire_2219});
or_n #(2, 0, 0) OR_317 (c6288_wire_1093, {c6288_wire_304, c6288_wire_2221});
nand_n #(2, 0, 0) NAND_67 (c6288_wire_2222, {c6288_wire_25_34, c6288_wire_114_36});
notg #(0, 0) NOT_329 (c6288_wire_2223, c6288_wire_305_1);
and_n #(2, 0, 0) AND_869 (c6288_wire_2221, {c6288_wire_2223, c6288_wire_2222});
or_n #(2, 0, 0) OR_318 (c6288_wire_1098, {c6288_wire_302, c6288_wire_2224});
nand_n #(2, 0, 0) NAND_68 (c6288_wire_2225, {c6288_wire_25_35, c6288_wire_117_36});
notg #(0, 0) NOT_330 (c6288_wire_2226, c6288_wire_303_1);
and_n #(2, 0, 0) AND_870 (c6288_wire_2224, {c6288_wire_2226, c6288_wire_2225});
nor_n #(2, 0, 0) NOR_7 (c6288_wire_1981, {c6288_wire_1104_1, c6288_wire_1103_3});
or_n #(2, 0, 0) OR_319 (c6288_wire_1109, {c6288_wire_2227, c6288_wire_2228});
notg #(0, 0) NOT_331 (c6288_wire_2229, c6288_wire_740_2);
and_n #(2, 0, 0) AND_871 (c6288_wire_2227, {c6288_wire_2229, c6288_wire_2230_0});
and_n #(2, 0, 0) AND_872 (c6288_wire_2228, {c6288_wire_288, c6288_wire_2231});
notg #(0, 0) NOT_332 (c6288_wire_2231, c6288_wire_2230_1);
or_n #(2, 0, 0) OR_320 (c6288_wire_1116, {c6288_wire_326, c6288_wire_2232});
nand_n #(2, 0, 0) NAND_69 (c6288_wire_2233, {c6288_wire_25_36, c6288_wire_81_36});
notg #(0, 0) NOT_333 (c6288_wire_2234, c6288_wire_327_1);
and_n #(2, 0, 0) AND_873 (c6288_wire_2232, {c6288_wire_2234, c6288_wire_2233});
or_n #(2, 0, 0) OR_321 (c6288_wire_1121, {c6288_wire_324, c6288_wire_2235});
nand_n #(2, 0, 0) NAND_70 (c6288_wire_2236, {c6288_wire_25_37, c6288_wire_84_36});
notg #(0, 0) NOT_334 (c6288_wire_2237, c6288_wire_325_1);
and_n #(2, 0, 0) AND_874 (c6288_wire_2235, {c6288_wire_2237, c6288_wire_2236});
or_n #(2, 0, 0) OR_322 (c6288_wire_1126, {c6288_wire_322, c6288_wire_2238});
nand_n #(2, 0, 0) NAND_71 (c6288_wire_2239, {c6288_wire_25_38, c6288_wire_87_36});
notg #(0, 0) NOT_335 (c6288_wire_2240, c6288_wire_323_1);
and_n #(2, 0, 0) AND_875 (c6288_wire_2238, {c6288_wire_2240, c6288_wire_2239});
or_n #(2, 0, 0) OR_323 (c6288_wire_1131, {c6288_wire_320, c6288_wire_2241});
nand_n #(2, 0, 0) NAND_72 (c6288_wire_2242, {c6288_wire_25_39, c6288_wire_90_36});
notg #(0, 0) NOT_336 (c6288_wire_2243, c6288_wire_321_1);
and_n #(2, 0, 0) AND_876 (c6288_wire_2241, {c6288_wire_2243, c6288_wire_2242});
or_n #(2, 0, 0) OR_324 (c6288_wire_1136, {c6288_wire_318, c6288_wire_2244});
nand_n #(2, 0, 0) NAND_73 (c6288_wire_2245, {c6288_wire_25_40, c6288_wire_93_36});
notg #(0, 0) NOT_337 (c6288_wire_2246, c6288_wire_319_1);
and_n #(2, 0, 0) AND_877 (c6288_wire_2244, {c6288_wire_2246, c6288_wire_2245});
or_n #(2, 0, 0) OR_325 (c6288_wire_1141, {c6288_wire_316, c6288_wire_2247});
nand_n #(2, 0, 0) NAND_74 (c6288_wire_2248, {c6288_wire_25_41, c6288_wire_96_36});
notg #(0, 0) NOT_338 (c6288_wire_2249, c6288_wire_317_1);
and_n #(2, 0, 0) AND_878 (c6288_wire_2247, {c6288_wire_2249, c6288_wire_2248});
or_n #(2, 0, 0) OR_326 (c6288_wire_1146, {c6288_wire_314, c6288_wire_2250});
nand_n #(2, 0, 0) NAND_75 (c6288_wire_2251, {c6288_wire_25_42, c6288_wire_99_36});
notg #(0, 0) NOT_339 (c6288_wire_2252, c6288_wire_315_1);
and_n #(2, 0, 0) AND_879 (c6288_wire_2250, {c6288_wire_2252, c6288_wire_2251});
or_n #(2, 0, 0) OR_327 (c6288_wire_1080, {c6288_wire_312, c6288_wire_2253});
nand_n #(2, 0, 0) NAND_76 (c6288_wire_2254, {c6288_wire_25_43, c6288_wire_102_36});
notg #(0, 0) NOT_340 (c6288_wire_2255, c6288_wire_313_1);
and_n #(2, 0, 0) AND_880 (c6288_wire_2253, {c6288_wire_2255, c6288_wire_2254});
or_n #(2, 0, 0) OR_328 (c6288_wire_746, {c6288_wire_40, c6288_wire_2256});
nand_n #(2, 0, 0) NAND_77 (c6288_wire_2257, {c6288_wire_30_31, c6288_wire_6_38});
and_n #(2, 0, 0) AND_881 (c6288_wire_2256, {c6288_wire_39, c6288_wire_2257});
or_n #(2, 0, 0) OR_329 (c6288_wire_750, {c6288_wire_383, c6288_wire_2258});
nand_n #(2, 0, 0) NAND_78 (c6288_wire_2259, {c6288_wire_30_32, c6288_wire_105_37});
notg #(0, 0) NOT_341 (c6288_wire_2260, c6288_wire_384_1);
and_n #(2, 0, 0) AND_882 (c6288_wire_2258, {c6288_wire_2260, c6288_wire_2259});
or_n #(2, 0, 0) OR_330 (c6288_wire_759, {c6288_wire_381, c6288_wire_2261});
nand_n #(2, 0, 0) NAND_79 (c6288_wire_2262, {c6288_wire_30_33, c6288_wire_108_37});
notg #(0, 0) NOT_342 (c6288_wire_2263, c6288_wire_382_1);
and_n #(2, 0, 0) AND_883 (c6288_wire_2261, {c6288_wire_2263, c6288_wire_2262});
or_n #(2, 0, 0) OR_331 (c6288_wire_765, {c6288_wire_379, c6288_wire_2264});
nand_n #(2, 0, 0) NAND_80 (c6288_wire_2265, {c6288_wire_30_34, c6288_wire_111_37});
notg #(0, 0) NOT_343 (c6288_wire_2266, c6288_wire_380_1);
and_n #(2, 0, 0) AND_884 (c6288_wire_2264, {c6288_wire_2266, c6288_wire_2265});
or_n #(2, 0, 0) OR_332 (c6288_wire_771, {c6288_wire_377, c6288_wire_2267});
nand_n #(2, 0, 0) NAND_81 (c6288_wire_2268, {c6288_wire_30_35, c6288_wire_114_37});
notg #(0, 0) NOT_344 (c6288_wire_2269, c6288_wire_378_1);
and_n #(2, 0, 0) AND_885 (c6288_wire_2267, {c6288_wire_2269, c6288_wire_2268});
or_n #(2, 0, 0) OR_333 (c6288_wire_777, {c6288_wire_375, c6288_wire_2270});
nand_n #(2, 0, 0) NAND_82 (c6288_wire_2271, {c6288_wire_30_36, c6288_wire_117_37});
notg #(0, 0) NOT_345 (c6288_wire_2272, c6288_wire_376_1);
and_n #(2, 0, 0) AND_886 (c6288_wire_2270, {c6288_wire_2272, c6288_wire_2271});
or_n #(2, 0, 0) OR_334 (c6288_wire_786, {c6288_wire_401, c6288_wire_2273});
nand_n #(2, 0, 0) NAND_83 (c6288_wire_2274, {c6288_wire_30_37, c6288_wire_78_37});
notg #(0, 0) NOT_346 (c6288_wire_2275, c6288_wire_402_1);
and_n #(2, 0, 0) AND_887 (c6288_wire_2273, {c6288_wire_2275, c6288_wire_2274});
or_n #(2, 0, 0) OR_335 (c6288_wire_793, {c6288_wire_399, c6288_wire_2276});
nand_n #(2, 0, 0) NAND_84 (c6288_wire_2277, {c6288_wire_30_38, c6288_wire_81_37});
notg #(0, 0) NOT_347 (c6288_wire_2278, c6288_wire_400_1);
and_n #(2, 0, 0) AND_888 (c6288_wire_2276, {c6288_wire_2278, c6288_wire_2277});
or_n #(2, 0, 0) OR_336 (c6288_wire_799, {c6288_wire_397, c6288_wire_2279});
nand_n #(2, 0, 0) NAND_85 (c6288_wire_2280, {c6288_wire_30_39, c6288_wire_84_37});
notg #(0, 0) NOT_348 (c6288_wire_2281, c6288_wire_398_1);
and_n #(2, 0, 0) AND_889 (c6288_wire_2279, {c6288_wire_2281, c6288_wire_2280});
or_n #(2, 0, 0) OR_337 (c6288_wire_805, {c6288_wire_395, c6288_wire_2282});
nand_n #(2, 0, 0) NAND_86 (c6288_wire_2283, {c6288_wire_30_40, c6288_wire_87_37});
notg #(0, 0) NOT_349 (c6288_wire_2284, c6288_wire_396_1);
and_n #(2, 0, 0) AND_890 (c6288_wire_2282, {c6288_wire_2284, c6288_wire_2283});
or_n #(2, 0, 0) OR_338 (c6288_wire_811, {c6288_wire_393, c6288_wire_2285});
nand_n #(2, 0, 0) NAND_87 (c6288_wire_2286, {c6288_wire_30_41, c6288_wire_90_37});
notg #(0, 0) NOT_350 (c6288_wire_2287, c6288_wire_394_1);
and_n #(2, 0, 0) AND_891 (c6288_wire_2285, {c6288_wire_2287, c6288_wire_2286});
or_n #(2, 0, 0) OR_339 (c6288_wire_817, {c6288_wire_391, c6288_wire_2288});
nand_n #(2, 0, 0) NAND_88 (c6288_wire_2289, {c6288_wire_30_42, c6288_wire_93_37});
notg #(0, 0) NOT_351 (c6288_wire_2290, c6288_wire_392_1);
and_n #(2, 0, 0) AND_892 (c6288_wire_2288, {c6288_wire_2290, c6288_wire_2289});
or_n #(2, 0, 0) OR_340 (c6288_wire_823, {c6288_wire_389, c6288_wire_2291});
nand_n #(2, 0, 0) NAND_89 (c6288_wire_2292, {c6288_wire_30_43, c6288_wire_96_37});
notg #(0, 0) NOT_352 (c6288_wire_2293, c6288_wire_390_1);
and_n #(2, 0, 0) AND_893 (c6288_wire_2291, {c6288_wire_2293, c6288_wire_2292});
or_n #(2, 0, 0) OR_341 (c6288_wire_829, {c6288_wire_387, c6288_wire_2294});
nand_n #(2, 0, 0) NAND_90 (c6288_wire_2295, {c6288_wire_30_44, c6288_wire_99_37});
notg #(0, 0) NOT_353 (c6288_wire_2296, c6288_wire_388_1);
and_n #(2, 0, 0) AND_894 (c6288_wire_2294, {c6288_wire_2296, c6288_wire_2295});
or_n #(2, 0, 0) OR_342 (c6288_wire_755, {c6288_wire_385, c6288_wire_2297});
nand_n #(2, 0, 0) NAND_91 (c6288_wire_2298, {c6288_wire_30_45, c6288_wire_102_37});
notg #(0, 0) NOT_354 (c6288_wire_2299, c6288_wire_386_1);
and_n #(2, 0, 0) AND_895 (c6288_wire_2297, {c6288_wire_2299, c6288_wire_2298});
or_n #(2, 0, 0) OR_343 (c6288_wire_1234, {c6288_wire_45, c6288_wire_2300});
nand_n #(2, 0, 0) NAND_92 (c6288_wire_2301, {c6288_wire_37_31, c6288_wire_6_39});
and_n #(2, 0, 0) AND_896 (c6288_wire_2300, {c6288_wire_44, c6288_wire_2301});
or_n #(2, 0, 0) OR_344 (c6288_wire_1237, {c6288_wire_425, c6288_wire_2302});
nand_n #(2, 0, 0) NAND_93 (c6288_wire_2303, {c6288_wire_37_32, c6288_wire_105_38});
notg #(0, 0) NOT_355 (c6288_wire_2304, c6288_wire_426_1);
and_n #(2, 0, 0) AND_897 (c6288_wire_2302, {c6288_wire_2304, c6288_wire_2303});
or_n #(2, 0, 0) OR_345 (c6288_wire_1245, {c6288_wire_423, c6288_wire_2305});
nand_n #(2, 0, 0) NAND_94 (c6288_wire_2306, {c6288_wire_37_33, c6288_wire_108_38});
notg #(0, 0) NOT_356 (c6288_wire_2307, c6288_wire_424_1);
and_n #(2, 0, 0) AND_898 (c6288_wire_2305, {c6288_wire_2307, c6288_wire_2306});
or_n #(2, 0, 0) OR_346 (c6288_wire_1250, {c6288_wire_421, c6288_wire_2308});
nand_n #(2, 0, 0) NAND_95 (c6288_wire_2309, {c6288_wire_37_34, c6288_wire_111_38});
notg #(0, 0) NOT_357 (c6288_wire_2310, c6288_wire_422_1);
and_n #(2, 0, 0) AND_899 (c6288_wire_2308, {c6288_wire_2310, c6288_wire_2309});
or_n #(2, 0, 0) OR_347 (c6288_wire_1255, {c6288_wire_419, c6288_wire_2311});
nand_n #(2, 0, 0) NAND_96 (c6288_wire_2312, {c6288_wire_37_35, c6288_wire_114_38});
notg #(0, 0) NOT_358 (c6288_wire_2313, c6288_wire_420_1);
and_n #(2, 0, 0) AND_900 (c6288_wire_2311, {c6288_wire_2313, c6288_wire_2312});
or_n #(2, 0, 0) OR_348 (c6288_wire_1260, {c6288_wire_417, c6288_wire_2314});
nand_n #(2, 0, 0) NAND_97 (c6288_wire_2315, {c6288_wire_37_36, c6288_wire_117_38});
notg #(0, 0) NOT_359 (c6288_wire_2316, c6288_wire_418_1);
and_n #(2, 0, 0) AND_901 (c6288_wire_2314, {c6288_wire_2316, c6288_wire_2315});
nor_n #(2, 0, 0) NOR_8 (c6288_wire_1952, {c6288_wire_1266_2, c6288_wire_1265_2});
or_n #(2, 0, 0) OR_349 (c6288_wire_1270, {c6288_wire_443, c6288_wire_2317});
nand_n #(2, 0, 0) NAND_98 (c6288_wire_2318, {c6288_wire_37_37, c6288_wire_78_38});
notg #(0, 0) NOT_360 (c6288_wire_2319, c6288_wire_444_1);
and_n #(2, 0, 0) AND_902 (c6288_wire_2317, {c6288_wire_2319, c6288_wire_2318});
or_n #(2, 0, 0) OR_350 (c6288_wire_1276, {c6288_wire_441, c6288_wire_2320});
nand_n #(2, 0, 0) NAND_99 (c6288_wire_2321, {c6288_wire_37_38, c6288_wire_81_38});
notg #(0, 0) NOT_361 (c6288_wire_2322, c6288_wire_442_1);
and_n #(2, 0, 0) AND_903 (c6288_wire_2320, {c6288_wire_2322, c6288_wire_2321});
or_n #(2, 0, 0) OR_351 (c6288_wire_1281, {c6288_wire_439, c6288_wire_2323});
nand_n #(2, 0, 0) NAND_100 (c6288_wire_2324, {c6288_wire_37_39, c6288_wire_84_38});
notg #(0, 0) NOT_362 (c6288_wire_2325, c6288_wire_440_1);
and_n #(2, 0, 0) AND_904 (c6288_wire_2323, {c6288_wire_2325, c6288_wire_2324});
or_n #(2, 0, 0) OR_352 (c6288_wire_1286, {c6288_wire_437, c6288_wire_2326});
nand_n #(2, 0, 0) NAND_101 (c6288_wire_2327, {c6288_wire_37_40, c6288_wire_87_38});
notg #(0, 0) NOT_363 (c6288_wire_2328, c6288_wire_438_1);
and_n #(2, 0, 0) AND_905 (c6288_wire_2326, {c6288_wire_2328, c6288_wire_2327});
or_n #(2, 0, 0) OR_353 (c6288_wire_1291, {c6288_wire_435, c6288_wire_2329});
nand_n #(2, 0, 0) NAND_102 (c6288_wire_2330, {c6288_wire_37_41, c6288_wire_90_38});
notg #(0, 0) NOT_364 (c6288_wire_2331, c6288_wire_436_1);
and_n #(2, 0, 0) AND_906 (c6288_wire_2329, {c6288_wire_2331, c6288_wire_2330});
or_n #(2, 0, 0) OR_354 (c6288_wire_1296, {c6288_wire_433, c6288_wire_2332});
nand_n #(2, 0, 0) NAND_103 (c6288_wire_2333, {c6288_wire_37_42, c6288_wire_93_38});
notg #(0, 0) NOT_365 (c6288_wire_2334, c6288_wire_434_1);
and_n #(2, 0, 0) AND_907 (c6288_wire_2332, {c6288_wire_2334, c6288_wire_2333});
or_n #(2, 0, 0) OR_355 (c6288_wire_1301, {c6288_wire_431, c6288_wire_2335});
nand_n #(2, 0, 0) NAND_104 (c6288_wire_2336, {c6288_wire_37_43, c6288_wire_96_38});
notg #(0, 0) NOT_366 (c6288_wire_2337, c6288_wire_432_1);
and_n #(2, 0, 0) AND_908 (c6288_wire_2335, {c6288_wire_2337, c6288_wire_2336});
or_n #(2, 0, 0) OR_356 (c6288_wire_1306, {c6288_wire_429, c6288_wire_2338});
nand_n #(2, 0, 0) NAND_105 (c6288_wire_2339, {c6288_wire_37_44, c6288_wire_99_38});
notg #(0, 0) NOT_367 (c6288_wire_2340, c6288_wire_430_1);
and_n #(2, 0, 0) AND_909 (c6288_wire_2338, {c6288_wire_2340, c6288_wire_2339});
or_n #(2, 0, 0) OR_357 (c6288_wire_1242, {c6288_wire_427, c6288_wire_2341});
nand_n #(2, 0, 0) NAND_106 (c6288_wire_2342, {c6288_wire_37_45, c6288_wire_102_38});
notg #(0, 0) NOT_368 (c6288_wire_2343, c6288_wire_428_1);
and_n #(2, 0, 0) AND_910 (c6288_wire_2341, {c6288_wire_2343, c6288_wire_2342});
or_n #(2, 0, 0) OR_358 (c6288_wire_1313, {c6288_wire_50, c6288_wire_2344});
nand_n #(2, 0, 0) NAND_107 (c6288_wire_2345, {c6288_wire_42_31, c6288_wire_6_40});
and_n #(2, 0, 0) AND_911 (c6288_wire_2344, {c6288_wire_49, c6288_wire_2345});
or_n #(2, 0, 0) OR_359 (c6288_wire_1316, {c6288_wire_467, c6288_wire_2346});
nand_n #(2, 0, 0) NAND_108 (c6288_wire_2347, {c6288_wire_42_32, c6288_wire_105_39});
notg #(0, 0) NOT_369 (c6288_wire_2348, c6288_wire_468_1);
and_n #(2, 0, 0) AND_912 (c6288_wire_2346, {c6288_wire_2348, c6288_wire_2347});
or_n #(2, 0, 0) OR_360 (c6288_wire_1324, {c6288_wire_465, c6288_wire_2349});
nand_n #(2, 0, 0) NAND_109 (c6288_wire_2350, {c6288_wire_42_33, c6288_wire_108_39});
notg #(0, 0) NOT_370 (c6288_wire_2351, c6288_wire_466_1);
and_n #(2, 0, 0) AND_913 (c6288_wire_2349, {c6288_wire_2351, c6288_wire_2350});
or_n #(2, 0, 0) OR_361 (c6288_wire_1329, {c6288_wire_463, c6288_wire_2352});
nand_n #(2, 0, 0) NAND_110 (c6288_wire_2353, {c6288_wire_42_34, c6288_wire_111_39});
notg #(0, 0) NOT_371 (c6288_wire_2354, c6288_wire_464_1);
and_n #(2, 0, 0) AND_914 (c6288_wire_2352, {c6288_wire_2354, c6288_wire_2353});
or_n #(2, 0, 0) OR_362 (c6288_wire_1334, {c6288_wire_461, c6288_wire_2355});
nand_n #(2, 0, 0) NAND_111 (c6288_wire_2356, {c6288_wire_42_35, c6288_wire_114_39});
notg #(0, 0) NOT_372 (c6288_wire_2357, c6288_wire_462_1);
and_n #(2, 0, 0) AND_915 (c6288_wire_2355, {c6288_wire_2357, c6288_wire_2356});
or_n #(2, 0, 0) OR_363 (c6288_wire_1339, {c6288_wire_459, c6288_wire_2358});
nand_n #(2, 0, 0) NAND_112 (c6288_wire_2359, {c6288_wire_42_36, c6288_wire_117_39});
notg #(0, 0) NOT_373 (c6288_wire_2360, c6288_wire_460_1);
and_n #(2, 0, 0) AND_916 (c6288_wire_2358, {c6288_wire_2360, c6288_wire_2359});
nor_n #(2, 0, 0) NOR_9 (c6288_wire_1954, {c6288_wire_1345_2, c6288_wire_1344_2});
or_n #(2, 0, 0) OR_364 (c6288_wire_1348, {c6288_wire_485, c6288_wire_2361});
nand_n #(2, 0, 0) NAND_113 (c6288_wire_2362, {c6288_wire_42_37, c6288_wire_78_39});
notg #(0, 0) NOT_374 (c6288_wire_2363, c6288_wire_486_1);
and_n #(2, 0, 0) AND_917 (c6288_wire_2361, {c6288_wire_2363, c6288_wire_2362});
or_n #(2, 0, 0) OR_365 (c6288_wire_1354, {c6288_wire_483, c6288_wire_2364});
nand_n #(2, 0, 0) NAND_114 (c6288_wire_2365, {c6288_wire_42_38, c6288_wire_81_39});
notg #(0, 0) NOT_375 (c6288_wire_2366, c6288_wire_484_1);
and_n #(2, 0, 0) AND_918 (c6288_wire_2364, {c6288_wire_2366, c6288_wire_2365});
or_n #(2, 0, 0) OR_366 (c6288_wire_1359, {c6288_wire_481, c6288_wire_2367});
nand_n #(2, 0, 0) NAND_115 (c6288_wire_2368, {c6288_wire_42_39, c6288_wire_84_39});
notg #(0, 0) NOT_376 (c6288_wire_2369, c6288_wire_482_1);
and_n #(2, 0, 0) AND_919 (c6288_wire_2367, {c6288_wire_2369, c6288_wire_2368});
or_n #(2, 0, 0) OR_367 (c6288_wire_1364, {c6288_wire_479, c6288_wire_2370});
nand_n #(2, 0, 0) NAND_116 (c6288_wire_2371, {c6288_wire_42_40, c6288_wire_87_39});
notg #(0, 0) NOT_377 (c6288_wire_2372, c6288_wire_480_1);
and_n #(2, 0, 0) AND_920 (c6288_wire_2370, {c6288_wire_2372, c6288_wire_2371});
or_n #(2, 0, 0) OR_368 (c6288_wire_1369, {c6288_wire_477, c6288_wire_2373});
nand_n #(2, 0, 0) NAND_117 (c6288_wire_2374, {c6288_wire_42_41, c6288_wire_90_39});
notg #(0, 0) NOT_378 (c6288_wire_2375, c6288_wire_478_1);
and_n #(2, 0, 0) AND_921 (c6288_wire_2373, {c6288_wire_2375, c6288_wire_2374});
or_n #(2, 0, 0) OR_369 (c6288_wire_1374, {c6288_wire_475, c6288_wire_2376});
nand_n #(2, 0, 0) NAND_118 (c6288_wire_2377, {c6288_wire_42_42, c6288_wire_93_39});
notg #(0, 0) NOT_379 (c6288_wire_2378, c6288_wire_476_1);
and_n #(2, 0, 0) AND_922 (c6288_wire_2376, {c6288_wire_2378, c6288_wire_2377});
or_n #(2, 0, 0) OR_370 (c6288_wire_1379, {c6288_wire_473, c6288_wire_2379});
nand_n #(2, 0, 0) NAND_119 (c6288_wire_2380, {c6288_wire_42_43, c6288_wire_96_39});
notg #(0, 0) NOT_380 (c6288_wire_2381, c6288_wire_474_1);
and_n #(2, 0, 0) AND_923 (c6288_wire_2379, {c6288_wire_2381, c6288_wire_2380});
or_n #(2, 0, 0) OR_371 (c6288_wire_1384, {c6288_wire_471, c6288_wire_2382});
nand_n #(2, 0, 0) NAND_120 (c6288_wire_2383, {c6288_wire_42_44, c6288_wire_99_39});
notg #(0, 0) NOT_381 (c6288_wire_2384, c6288_wire_472_1);
and_n #(2, 0, 0) AND_924 (c6288_wire_2382, {c6288_wire_2384, c6288_wire_2383});
or_n #(2, 0, 0) OR_372 (c6288_wire_1321, {c6288_wire_469, c6288_wire_2385});
nand_n #(2, 0, 0) NAND_121 (c6288_wire_2386, {c6288_wire_42_45, c6288_wire_102_39});
notg #(0, 0) NOT_382 (c6288_wire_2387, c6288_wire_470_1);
and_n #(2, 0, 0) AND_925 (c6288_wire_2385, {c6288_wire_2387, c6288_wire_2386});
or_n #(2, 0, 0) OR_373 (c6288_wire_1391, {c6288_wire_55, c6288_wire_2388});
nand_n #(2, 0, 0) NAND_122 (c6288_wire_2389, {c6288_wire_47_31, c6288_wire_6_41});
and_n #(2, 0, 0) AND_926 (c6288_wire_2388, {c6288_wire_54, c6288_wire_2389});
or_n #(2, 0, 0) OR_374 (c6288_wire_1394, {c6288_wire_509, c6288_wire_2390});
nand_n #(2, 0, 0) NAND_123 (c6288_wire_2391, {c6288_wire_47_32, c6288_wire_105_40});
notg #(0, 0) NOT_383 (c6288_wire_2392, c6288_wire_510_1);
and_n #(2, 0, 0) AND_927 (c6288_wire_2390, {c6288_wire_2392, c6288_wire_2391});
or_n #(2, 0, 0) OR_375 (c6288_wire_1402, {c6288_wire_507, c6288_wire_2393});
nand_n #(2, 0, 0) NAND_124 (c6288_wire_2394, {c6288_wire_47_33, c6288_wire_108_40});
notg #(0, 0) NOT_384 (c6288_wire_2395, c6288_wire_508_1);
and_n #(2, 0, 0) AND_928 (c6288_wire_2393, {c6288_wire_2395, c6288_wire_2394});
or_n #(2, 0, 0) OR_376 (c6288_wire_1407, {c6288_wire_505, c6288_wire_2396});
nand_n #(2, 0, 0) NAND_125 (c6288_wire_2397, {c6288_wire_47_34, c6288_wire_111_40});
notg #(0, 0) NOT_385 (c6288_wire_2398, c6288_wire_506_1);
and_n #(2, 0, 0) AND_929 (c6288_wire_2396, {c6288_wire_2398, c6288_wire_2397});
or_n #(2, 0, 0) OR_377 (c6288_wire_1412, {c6288_wire_503, c6288_wire_2399});
nand_n #(2, 0, 0) NAND_126 (c6288_wire_2400, {c6288_wire_47_35, c6288_wire_114_40});
notg #(0, 0) NOT_386 (c6288_wire_2401, c6288_wire_504_1);
and_n #(2, 0, 0) AND_930 (c6288_wire_2399, {c6288_wire_2401, c6288_wire_2400});
or_n #(2, 0, 0) OR_378 (c6288_wire_1417, {c6288_wire_501, c6288_wire_2402});
nand_n #(2, 0, 0) NAND_127 (c6288_wire_2403, {c6288_wire_47_36, c6288_wire_117_40});
notg #(0, 0) NOT_387 (c6288_wire_2404, c6288_wire_502_1);
and_n #(2, 0, 0) AND_931 (c6288_wire_2402, {c6288_wire_2404, c6288_wire_2403});
nor_n #(2, 0, 0) NOR_10 (c6288_wire_1958, {c6288_wire_1423_2, c6288_wire_1422_2});
or_n #(2, 0, 0) OR_379 (c6288_wire_1426, {c6288_wire_527, c6288_wire_2405});
nand_n #(2, 0, 0) NAND_128 (c6288_wire_2406, {c6288_wire_47_37, c6288_wire_78_40});
notg #(0, 0) NOT_388 (c6288_wire_2407, c6288_wire_528_1);
and_n #(2, 0, 0) AND_932 (c6288_wire_2405, {c6288_wire_2407, c6288_wire_2406});
or_n #(2, 0, 0) OR_380 (c6288_wire_1432, {c6288_wire_525, c6288_wire_2408});
nand_n #(2, 0, 0) NAND_129 (c6288_wire_2409, {c6288_wire_47_38, c6288_wire_81_40});
notg #(0, 0) NOT_389 (c6288_wire_2410, c6288_wire_526_1);
and_n #(2, 0, 0) AND_933 (c6288_wire_2408, {c6288_wire_2410, c6288_wire_2409});
or_n #(2, 0, 0) OR_381 (c6288_wire_1437, {c6288_wire_523, c6288_wire_2411});
nand_n #(2, 0, 0) NAND_130 (c6288_wire_2412, {c6288_wire_47_39, c6288_wire_84_40});
notg #(0, 0) NOT_390 (c6288_wire_2413, c6288_wire_524_1);
and_n #(2, 0, 0) AND_934 (c6288_wire_2411, {c6288_wire_2413, c6288_wire_2412});
or_n #(2, 0, 0) OR_382 (c6288_wire_1442, {c6288_wire_521, c6288_wire_2414});
nand_n #(2, 0, 0) NAND_131 (c6288_wire_2415, {c6288_wire_47_40, c6288_wire_87_40});
notg #(0, 0) NOT_391 (c6288_wire_2416, c6288_wire_522_1);
and_n #(2, 0, 0) AND_935 (c6288_wire_2414, {c6288_wire_2416, c6288_wire_2415});
or_n #(2, 0, 0) OR_383 (c6288_wire_1447, {c6288_wire_519, c6288_wire_2417});
nand_n #(2, 0, 0) NAND_132 (c6288_wire_2418, {c6288_wire_47_41, c6288_wire_90_40});
notg #(0, 0) NOT_392 (c6288_wire_2419, c6288_wire_520_1);
and_n #(2, 0, 0) AND_936 (c6288_wire_2417, {c6288_wire_2419, c6288_wire_2418});
or_n #(2, 0, 0) OR_384 (c6288_wire_1452, {c6288_wire_517, c6288_wire_2420});
nand_n #(2, 0, 0) NAND_133 (c6288_wire_2421, {c6288_wire_47_42, c6288_wire_93_40});
notg #(0, 0) NOT_393 (c6288_wire_2422, c6288_wire_518_1);
and_n #(2, 0, 0) AND_937 (c6288_wire_2420, {c6288_wire_2422, c6288_wire_2421});
or_n #(2, 0, 0) OR_385 (c6288_wire_1457, {c6288_wire_515, c6288_wire_2423});
nand_n #(2, 0, 0) NAND_134 (c6288_wire_2424, {c6288_wire_47_43, c6288_wire_96_40});
notg #(0, 0) NOT_394 (c6288_wire_2425, c6288_wire_516_1);
and_n #(2, 0, 0) AND_938 (c6288_wire_2423, {c6288_wire_2425, c6288_wire_2424});
or_n #(2, 0, 0) OR_386 (c6288_wire_1462, {c6288_wire_513, c6288_wire_2426});
nand_n #(2, 0, 0) NAND_135 (c6288_wire_2427, {c6288_wire_47_44, c6288_wire_99_40});
notg #(0, 0) NOT_395 (c6288_wire_2428, c6288_wire_514_1);
and_n #(2, 0, 0) AND_939 (c6288_wire_2426, {c6288_wire_2428, c6288_wire_2427});
or_n #(2, 0, 0) OR_387 (c6288_wire_1399, {c6288_wire_511, c6288_wire_2429});
nand_n #(2, 0, 0) NAND_136 (c6288_wire_2430, {c6288_wire_47_45, c6288_wire_102_40});
notg #(0, 0) NOT_396 (c6288_wire_2431, c6288_wire_512_1);
and_n #(2, 0, 0) AND_940 (c6288_wire_2429, {c6288_wire_2431, c6288_wire_2430});
or_n #(2, 0, 0) OR_388 (c6288_wire_1469, {c6288_wire_60, c6288_wire_2432});
nand_n #(2, 0, 0) NAND_137 (c6288_wire_2433, {c6288_wire_52_31, c6288_wire_6_42});
and_n #(2, 0, 0) AND_941 (c6288_wire_2432, {c6288_wire_59, c6288_wire_2433});
or_n #(2, 0, 0) OR_389 (c6288_wire_1472, {c6288_wire_551, c6288_wire_2434});
nand_n #(2, 0, 0) NAND_138 (c6288_wire_2435, {c6288_wire_52_32, c6288_wire_105_41});
notg #(0, 0) NOT_397 (c6288_wire_2436, c6288_wire_552_1);
and_n #(2, 0, 0) AND_942 (c6288_wire_2434, {c6288_wire_2436, c6288_wire_2435});
or_n #(2, 0, 0) OR_390 (c6288_wire_1480, {c6288_wire_549, c6288_wire_2437});
nand_n #(2, 0, 0) NAND_139 (c6288_wire_2438, {c6288_wire_52_33, c6288_wire_108_41});
notg #(0, 0) NOT_398 (c6288_wire_2439, c6288_wire_550_1);
and_n #(2, 0, 0) AND_943 (c6288_wire_2437, {c6288_wire_2439, c6288_wire_2438});
or_n #(2, 0, 0) OR_391 (c6288_wire_1485, {c6288_wire_547, c6288_wire_2440});
nand_n #(2, 0, 0) NAND_140 (c6288_wire_2441, {c6288_wire_52_34, c6288_wire_111_41});
notg #(0, 0) NOT_399 (c6288_wire_2442, c6288_wire_548_1);
and_n #(2, 0, 0) AND_944 (c6288_wire_2440, {c6288_wire_2442, c6288_wire_2441});
or_n #(2, 0, 0) OR_392 (c6288_wire_1490, {c6288_wire_545, c6288_wire_2443});
nand_n #(2, 0, 0) NAND_141 (c6288_wire_2444, {c6288_wire_52_35, c6288_wire_114_41});
notg #(0, 0) NOT_400 (c6288_wire_2445, c6288_wire_546_1);
and_n #(2, 0, 0) AND_945 (c6288_wire_2443, {c6288_wire_2445, c6288_wire_2444});
or_n #(2, 0, 0) OR_393 (c6288_wire_1495, {c6288_wire_543, c6288_wire_2446});
nand_n #(2, 0, 0) NAND_142 (c6288_wire_2447, {c6288_wire_52_36, c6288_wire_117_41});
notg #(0, 0) NOT_401 (c6288_wire_2448, c6288_wire_544_1);
and_n #(2, 0, 0) AND_946 (c6288_wire_2446, {c6288_wire_2448, c6288_wire_2447});
nor_n #(2, 0, 0) NOR_11 (c6288_wire_1960, {c6288_wire_1501_2, c6288_wire_1500_2});
or_n #(2, 0, 0) OR_394 (c6288_wire_1504, {c6288_wire_569, c6288_wire_2449});
nand_n #(2, 0, 0) NAND_143 (c6288_wire_2450, {c6288_wire_52_37, c6288_wire_78_41});
notg #(0, 0) NOT_402 (c6288_wire_2451, c6288_wire_570_1);
and_n #(2, 0, 0) AND_947 (c6288_wire_2449, {c6288_wire_2451, c6288_wire_2450});
or_n #(2, 0, 0) OR_395 (c6288_wire_1510, {c6288_wire_567, c6288_wire_2452});
nand_n #(2, 0, 0) NAND_144 (c6288_wire_2453, {c6288_wire_52_38, c6288_wire_81_41});
notg #(0, 0) NOT_403 (c6288_wire_2454, c6288_wire_568_1);
and_n #(2, 0, 0) AND_948 (c6288_wire_2452, {c6288_wire_2454, c6288_wire_2453});
or_n #(2, 0, 0) OR_396 (c6288_wire_1515, {c6288_wire_565, c6288_wire_2455});
nand_n #(2, 0, 0) NAND_145 (c6288_wire_2456, {c6288_wire_52_39, c6288_wire_84_41});
notg #(0, 0) NOT_404 (c6288_wire_2457, c6288_wire_566_1);
and_n #(2, 0, 0) AND_949 (c6288_wire_2455, {c6288_wire_2457, c6288_wire_2456});
or_n #(2, 0, 0) OR_397 (c6288_wire_1520, {c6288_wire_563, c6288_wire_2458});
nand_n #(2, 0, 0) NAND_146 (c6288_wire_2459, {c6288_wire_52_40, c6288_wire_87_41});
notg #(0, 0) NOT_405 (c6288_wire_2460, c6288_wire_564_1);
and_n #(2, 0, 0) AND_950 (c6288_wire_2458, {c6288_wire_2460, c6288_wire_2459});
or_n #(2, 0, 0) OR_398 (c6288_wire_1525, {c6288_wire_561, c6288_wire_2461});
nand_n #(2, 0, 0) NAND_147 (c6288_wire_2462, {c6288_wire_52_41, c6288_wire_90_41});
notg #(0, 0) NOT_406 (c6288_wire_2463, c6288_wire_562_1);
and_n #(2, 0, 0) AND_951 (c6288_wire_2461, {c6288_wire_2463, c6288_wire_2462});
or_n #(2, 0, 0) OR_399 (c6288_wire_1530, {c6288_wire_559, c6288_wire_2464});
nand_n #(2, 0, 0) NAND_148 (c6288_wire_2465, {c6288_wire_52_42, c6288_wire_93_41});
notg #(0, 0) NOT_407 (c6288_wire_2466, c6288_wire_560_1);
and_n #(2, 0, 0) AND_952 (c6288_wire_2464, {c6288_wire_2466, c6288_wire_2465});
or_n #(2, 0, 0) OR_400 (c6288_wire_1535, {c6288_wire_557, c6288_wire_2467});
nand_n #(2, 0, 0) NAND_149 (c6288_wire_2468, {c6288_wire_52_43, c6288_wire_96_41});
notg #(0, 0) NOT_408 (c6288_wire_2469, c6288_wire_558_1);
and_n #(2, 0, 0) AND_953 (c6288_wire_2467, {c6288_wire_2469, c6288_wire_2468});
or_n #(2, 0, 0) OR_401 (c6288_wire_1540, {c6288_wire_555, c6288_wire_2470});
nand_n #(2, 0, 0) NAND_150 (c6288_wire_2471, {c6288_wire_52_44, c6288_wire_99_41});
notg #(0, 0) NOT_409 (c6288_wire_2472, c6288_wire_556_1);
and_n #(2, 0, 0) AND_954 (c6288_wire_2470, {c6288_wire_2472, c6288_wire_2471});
or_n #(2, 0, 0) OR_402 (c6288_wire_1477, {c6288_wire_553, c6288_wire_2473});
nand_n #(2, 0, 0) NAND_151 (c6288_wire_2474, {c6288_wire_52_45, c6288_wire_102_41});
notg #(0, 0) NOT_410 (c6288_wire_2475, c6288_wire_554_1);
and_n #(2, 0, 0) AND_955 (c6288_wire_2473, {c6288_wire_2475, c6288_wire_2474});
or_n #(2, 0, 0) OR_403 (c6288_wire_1547, {c6288_wire_65, c6288_wire_2476});
nand_n #(2, 0, 0) NAND_152 (c6288_wire_2477, {c6288_wire_57_31, c6288_wire_6_43});
and_n #(2, 0, 0) AND_956 (c6288_wire_2476, {c6288_wire_64, c6288_wire_2477});
or_n #(2, 0, 0) OR_404 (c6288_wire_1550, {c6288_wire_593, c6288_wire_2478});
nand_n #(2, 0, 0) NAND_153 (c6288_wire_2479, {c6288_wire_57_32, c6288_wire_105_42});
notg #(0, 0) NOT_411 (c6288_wire_2480, c6288_wire_594_1);
and_n #(2, 0, 0) AND_957 (c6288_wire_2478, {c6288_wire_2480, c6288_wire_2479});
or_n #(2, 0, 0) OR_405 (c6288_wire_1558, {c6288_wire_591, c6288_wire_2481});
nand_n #(2, 0, 0) NAND_154 (c6288_wire_2482, {c6288_wire_57_33, c6288_wire_108_42});
notg #(0, 0) NOT_412 (c6288_wire_2483, c6288_wire_592_1);
and_n #(2, 0, 0) AND_958 (c6288_wire_2481, {c6288_wire_2483, c6288_wire_2482});
or_n #(2, 0, 0) OR_406 (c6288_wire_1563, {c6288_wire_589, c6288_wire_2484});
nand_n #(2, 0, 0) NAND_155 (c6288_wire_2485, {c6288_wire_57_34, c6288_wire_111_42});
notg #(0, 0) NOT_413 (c6288_wire_2486, c6288_wire_590_1);
and_n #(2, 0, 0) AND_959 (c6288_wire_2484, {c6288_wire_2486, c6288_wire_2485});
or_n #(2, 0, 0) OR_407 (c6288_wire_1568, {c6288_wire_587, c6288_wire_2487});
nand_n #(2, 0, 0) NAND_156 (c6288_wire_2488, {c6288_wire_57_35, c6288_wire_114_42});
notg #(0, 0) NOT_414 (c6288_wire_2489, c6288_wire_588_1);
and_n #(2, 0, 0) AND_960 (c6288_wire_2487, {c6288_wire_2489, c6288_wire_2488});
or_n #(2, 0, 0) OR_408 (c6288_wire_1573, {c6288_wire_585, c6288_wire_2490});
nand_n #(2, 0, 0) NAND_157 (c6288_wire_2491, {c6288_wire_57_36, c6288_wire_117_42});
notg #(0, 0) NOT_415 (c6288_wire_2492, c6288_wire_586_1);
and_n #(2, 0, 0) AND_961 (c6288_wire_2490, {c6288_wire_2492, c6288_wire_2491});
nor_n #(2, 0, 0) NOR_12 (c6288_wire_1962, {c6288_wire_1579_2, c6288_wire_1578_2});
or_n #(2, 0, 0) OR_409 (c6288_wire_1582, {c6288_wire_611, c6288_wire_2493});
nand_n #(2, 0, 0) NAND_158 (c6288_wire_2494, {c6288_wire_57_37, c6288_wire_78_42});
notg #(0, 0) NOT_416 (c6288_wire_2495, c6288_wire_612_1);
and_n #(2, 0, 0) AND_962 (c6288_wire_2493, {c6288_wire_2495, c6288_wire_2494});
or_n #(2, 0, 0) OR_410 (c6288_wire_1588, {c6288_wire_609, c6288_wire_2496});
nand_n #(2, 0, 0) NAND_159 (c6288_wire_2497, {c6288_wire_57_38, c6288_wire_81_42});
notg #(0, 0) NOT_417 (c6288_wire_2498, c6288_wire_610_1);
and_n #(2, 0, 0) AND_963 (c6288_wire_2496, {c6288_wire_2498, c6288_wire_2497});
or_n #(2, 0, 0) OR_411 (c6288_wire_1593, {c6288_wire_607, c6288_wire_2499});
nand_n #(2, 0, 0) NAND_160 (c6288_wire_2500, {c6288_wire_57_39, c6288_wire_84_42});
notg #(0, 0) NOT_418 (c6288_wire_2501, c6288_wire_608_1);
and_n #(2, 0, 0) AND_964 (c6288_wire_2499, {c6288_wire_2501, c6288_wire_2500});
or_n #(2, 0, 0) OR_412 (c6288_wire_1598, {c6288_wire_605, c6288_wire_2502});
nand_n #(2, 0, 0) NAND_161 (c6288_wire_2503, {c6288_wire_57_40, c6288_wire_87_42});
notg #(0, 0) NOT_419 (c6288_wire_2504, c6288_wire_606_1);
and_n #(2, 0, 0) AND_965 (c6288_wire_2502, {c6288_wire_2504, c6288_wire_2503});
or_n #(2, 0, 0) OR_413 (c6288_wire_1603, {c6288_wire_603, c6288_wire_2505});
nand_n #(2, 0, 0) NAND_162 (c6288_wire_2506, {c6288_wire_57_41, c6288_wire_90_42});
notg #(0, 0) NOT_420 (c6288_wire_2507, c6288_wire_604_1);
and_n #(2, 0, 0) AND_966 (c6288_wire_2505, {c6288_wire_2507, c6288_wire_2506});
or_n #(2, 0, 0) OR_414 (c6288_wire_1608, {c6288_wire_601, c6288_wire_2508});
nand_n #(2, 0, 0) NAND_163 (c6288_wire_2509, {c6288_wire_57_42, c6288_wire_93_42});
notg #(0, 0) NOT_421 (c6288_wire_2510, c6288_wire_602_1);
and_n #(2, 0, 0) AND_967 (c6288_wire_2508, {c6288_wire_2510, c6288_wire_2509});
or_n #(2, 0, 0) OR_415 (c6288_wire_1613, {c6288_wire_599, c6288_wire_2511});
nand_n #(2, 0, 0) NAND_164 (c6288_wire_2512, {c6288_wire_57_43, c6288_wire_96_42});
notg #(0, 0) NOT_422 (c6288_wire_2513, c6288_wire_600_1);
and_n #(2, 0, 0) AND_968 (c6288_wire_2511, {c6288_wire_2513, c6288_wire_2512});
or_n #(2, 0, 0) OR_416 (c6288_wire_1618, {c6288_wire_597, c6288_wire_2514});
nand_n #(2, 0, 0) NAND_165 (c6288_wire_2515, {c6288_wire_57_44, c6288_wire_99_42});
notg #(0, 0) NOT_423 (c6288_wire_2516, c6288_wire_598_1);
and_n #(2, 0, 0) AND_969 (c6288_wire_2514, {c6288_wire_2516, c6288_wire_2515});
or_n #(2, 0, 0) OR_417 (c6288_wire_1555, {c6288_wire_595, c6288_wire_2517});
nand_n #(2, 0, 0) NAND_166 (c6288_wire_2518, {c6288_wire_57_45, c6288_wire_102_42});
notg #(0, 0) NOT_424 (c6288_wire_2519, c6288_wire_596_1);
and_n #(2, 0, 0) AND_970 (c6288_wire_2517, {c6288_wire_2519, c6288_wire_2518});
or_n #(2, 0, 0) OR_418 (c6288_wire_1625, {c6288_wire_70, c6288_wire_2520});
nand_n #(2, 0, 0) NAND_167 (c6288_wire_2521, {c6288_wire_62_31, c6288_wire_6_44});
and_n #(2, 0, 0) AND_971 (c6288_wire_2520, {c6288_wire_69, c6288_wire_2521});
or_n #(2, 0, 0) OR_419 (c6288_wire_1628, {c6288_wire_635, c6288_wire_2522});
nand_n #(2, 0, 0) NAND_168 (c6288_wire_2523, {c6288_wire_62_32, c6288_wire_105_43});
notg #(0, 0) NOT_425 (c6288_wire_2524, c6288_wire_636_1);
and_n #(2, 0, 0) AND_972 (c6288_wire_2522, {c6288_wire_2524, c6288_wire_2523});
or_n #(2, 0, 0) OR_420 (c6288_wire_1636, {c6288_wire_633, c6288_wire_2525});
nand_n #(2, 0, 0) NAND_169 (c6288_wire_2526, {c6288_wire_62_33, c6288_wire_108_43});
notg #(0, 0) NOT_426 (c6288_wire_2527, c6288_wire_634_1);
and_n #(2, 0, 0) AND_973 (c6288_wire_2525, {c6288_wire_2527, c6288_wire_2526});
or_n #(2, 0, 0) OR_421 (c6288_wire_1641, {c6288_wire_631, c6288_wire_2528});
nand_n #(2, 0, 0) NAND_170 (c6288_wire_2529, {c6288_wire_62_34, c6288_wire_111_43});
notg #(0, 0) NOT_427 (c6288_wire_2530, c6288_wire_632_1);
and_n #(2, 0, 0) AND_974 (c6288_wire_2528, {c6288_wire_2530, c6288_wire_2529});
or_n #(2, 0, 0) OR_422 (c6288_wire_1646, {c6288_wire_629, c6288_wire_2531});
nand_n #(2, 0, 0) NAND_171 (c6288_wire_2532, {c6288_wire_62_35, c6288_wire_114_43});
notg #(0, 0) NOT_428 (c6288_wire_2533, c6288_wire_630_1);
and_n #(2, 0, 0) AND_975 (c6288_wire_2531, {c6288_wire_2533, c6288_wire_2532});
or_n #(2, 0, 0) OR_423 (c6288_wire_1651, {c6288_wire_627, c6288_wire_2534});
nand_n #(2, 0, 0) NAND_172 (c6288_wire_2535, {c6288_wire_62_36, c6288_wire_117_43});
notg #(0, 0) NOT_429 (c6288_wire_2536, c6288_wire_628_1);
and_n #(2, 0, 0) AND_976 (c6288_wire_2534, {c6288_wire_2536, c6288_wire_2535});
nor_n #(2, 0, 0) NOR_13 (c6288_wire_1964, {c6288_wire_1657_2, c6288_wire_1656_2});
or_n #(2, 0, 0) OR_424 (c6288_wire_1660, {c6288_wire_653, c6288_wire_2537});
nand_n #(2, 0, 0) NAND_173 (c6288_wire_2538, {c6288_wire_62_37, c6288_wire_78_43});
notg #(0, 0) NOT_430 (c6288_wire_2539, c6288_wire_654_1);
and_n #(2, 0, 0) AND_977 (c6288_wire_2537, {c6288_wire_2539, c6288_wire_2538});
or_n #(2, 0, 0) OR_425 (c6288_wire_1666, {c6288_wire_651, c6288_wire_2540});
nand_n #(2, 0, 0) NAND_174 (c6288_wire_2541, {c6288_wire_62_38, c6288_wire_81_43});
notg #(0, 0) NOT_431 (c6288_wire_2542, c6288_wire_652_1);
and_n #(2, 0, 0) AND_978 (c6288_wire_2540, {c6288_wire_2542, c6288_wire_2541});
or_n #(2, 0, 0) OR_426 (c6288_wire_1671, {c6288_wire_649, c6288_wire_2543});
nand_n #(2, 0, 0) NAND_175 (c6288_wire_2544, {c6288_wire_62_39, c6288_wire_84_43});
notg #(0, 0) NOT_432 (c6288_wire_2545, c6288_wire_650_1);
and_n #(2, 0, 0) AND_979 (c6288_wire_2543, {c6288_wire_2545, c6288_wire_2544});
or_n #(2, 0, 0) OR_427 (c6288_wire_1676, {c6288_wire_647, c6288_wire_2546});
nand_n #(2, 0, 0) NAND_176 (c6288_wire_2547, {c6288_wire_62_40, c6288_wire_87_43});
notg #(0, 0) NOT_433 (c6288_wire_2548, c6288_wire_648_1);
and_n #(2, 0, 0) AND_980 (c6288_wire_2546, {c6288_wire_2548, c6288_wire_2547});
or_n #(2, 0, 0) OR_428 (c6288_wire_1681, {c6288_wire_645, c6288_wire_2549});
nand_n #(2, 0, 0) NAND_177 (c6288_wire_2550, {c6288_wire_62_41, c6288_wire_90_43});
notg #(0, 0) NOT_434 (c6288_wire_2551, c6288_wire_646_1);
and_n #(2, 0, 0) AND_981 (c6288_wire_2549, {c6288_wire_2551, c6288_wire_2550});
or_n #(2, 0, 0) OR_429 (c6288_wire_1686, {c6288_wire_643, c6288_wire_2552});
nand_n #(2, 0, 0) NAND_178 (c6288_wire_2553, {c6288_wire_62_42, c6288_wire_93_43});
notg #(0, 0) NOT_435 (c6288_wire_2554, c6288_wire_644_1);
and_n #(2, 0, 0) AND_982 (c6288_wire_2552, {c6288_wire_2554, c6288_wire_2553});
or_n #(2, 0, 0) OR_430 (c6288_wire_1691, {c6288_wire_641, c6288_wire_2555});
nand_n #(2, 0, 0) NAND_179 (c6288_wire_2556, {c6288_wire_62_43, c6288_wire_96_43});
notg #(0, 0) NOT_436 (c6288_wire_2557, c6288_wire_642_1);
and_n #(2, 0, 0) AND_983 (c6288_wire_2555, {c6288_wire_2557, c6288_wire_2556});
or_n #(2, 0, 0) OR_431 (c6288_wire_1696, {c6288_wire_639, c6288_wire_2558});
nand_n #(2, 0, 0) NAND_180 (c6288_wire_2559, {c6288_wire_62_44, c6288_wire_99_43});
notg #(0, 0) NOT_437 (c6288_wire_2560, c6288_wire_640_1);
and_n #(2, 0, 0) AND_984 (c6288_wire_2558, {c6288_wire_2560, c6288_wire_2559});
or_n #(2, 0, 0) OR_432 (c6288_wire_1633, {c6288_wire_637, c6288_wire_2561});
nand_n #(2, 0, 0) NAND_181 (c6288_wire_2562, {c6288_wire_62_45, c6288_wire_102_43});
notg #(0, 0) NOT_438 (c6288_wire_2563, c6288_wire_638_1);
and_n #(2, 0, 0) AND_985 (c6288_wire_2561, {c6288_wire_2563, c6288_wire_2562});
or_n #(2, 0, 0) OR_433 (c6288_wire_1703, {c6288_wire_74, c6288_wire_2564});
nand_n #(2, 0, 0) NAND_182 (c6288_wire_2565, {c6288_wire_67_31, c6288_wire_6_45});
and_n #(2, 0, 0) AND_986 (c6288_wire_2564, {c6288_wire_73, c6288_wire_2565});
or_n #(2, 0, 0) OR_434 (c6288_wire_1706, {c6288_wire_677, c6288_wire_2566});
nand_n #(2, 0, 0) NAND_183 (c6288_wire_2567, {c6288_wire_67_32, c6288_wire_105_44});
notg #(0, 0) NOT_439 (c6288_wire_2568, c6288_wire_678_1);
and_n #(2, 0, 0) AND_987 (c6288_wire_2566, {c6288_wire_2568, c6288_wire_2567});
or_n #(2, 0, 0) OR_435 (c6288_wire_1714, {c6288_wire_675, c6288_wire_2569});
nand_n #(2, 0, 0) NAND_184 (c6288_wire_2570, {c6288_wire_67_33, c6288_wire_108_44});
notg #(0, 0) NOT_440 (c6288_wire_2571, c6288_wire_676_1);
and_n #(2, 0, 0) AND_988 (c6288_wire_2569, {c6288_wire_2571, c6288_wire_2570});
or_n #(2, 0, 0) OR_436 (c6288_wire_1719, {c6288_wire_673, c6288_wire_2572});
nand_n #(2, 0, 0) NAND_185 (c6288_wire_2573, {c6288_wire_67_34, c6288_wire_111_44});
notg #(0, 0) NOT_441 (c6288_wire_2574, c6288_wire_674_1);
and_n #(2, 0, 0) AND_989 (c6288_wire_2572, {c6288_wire_2574, c6288_wire_2573});
or_n #(2, 0, 0) OR_437 (c6288_wire_1724, {c6288_wire_671, c6288_wire_2575});
nand_n #(2, 0, 0) NAND_186 (c6288_wire_2576, {c6288_wire_67_35, c6288_wire_114_44});
notg #(0, 0) NOT_442 (c6288_wire_2577, c6288_wire_672_1);
and_n #(2, 0, 0) AND_990 (c6288_wire_2575, {c6288_wire_2577, c6288_wire_2576});
or_n #(2, 0, 0) OR_438 (c6288_wire_1729, {c6288_wire_669, c6288_wire_2578});
nand_n #(2, 0, 0) NAND_187 (c6288_wire_2579, {c6288_wire_67_36, c6288_wire_117_44});
notg #(0, 0) NOT_443 (c6288_wire_2580, c6288_wire_670_1);
and_n #(2, 0, 0) AND_991 (c6288_wire_2578, {c6288_wire_2580, c6288_wire_2579});
nor_n #(2, 0, 0) NOR_14 (c6288_wire_1966, {c6288_wire_1735_2, c6288_wire_1734_2});
or_n #(2, 0, 0) OR_439 (c6288_wire_1738, {c6288_wire_695, c6288_wire_2581});
nand_n #(2, 0, 0) NAND_188 (c6288_wire_2582, {c6288_wire_67_37, c6288_wire_78_44});
notg #(0, 0) NOT_444 (c6288_wire_2583, c6288_wire_696_1);
and_n #(2, 0, 0) AND_992 (c6288_wire_2581, {c6288_wire_2583, c6288_wire_2582});
or_n #(2, 0, 0) OR_440 (c6288_wire_1744, {c6288_wire_693, c6288_wire_2584});
nand_n #(2, 0, 0) NAND_189 (c6288_wire_2585, {c6288_wire_67_38, c6288_wire_81_44});
notg #(0, 0) NOT_445 (c6288_wire_2586, c6288_wire_694_1);
and_n #(2, 0, 0) AND_993 (c6288_wire_2584, {c6288_wire_2586, c6288_wire_2585});
or_n #(2, 0, 0) OR_441 (c6288_wire_1749, {c6288_wire_691, c6288_wire_2587});
nand_n #(2, 0, 0) NAND_190 (c6288_wire_2588, {c6288_wire_67_39, c6288_wire_84_44});
notg #(0, 0) NOT_446 (c6288_wire_2589, c6288_wire_692_1);
and_n #(2, 0, 0) AND_994 (c6288_wire_2587, {c6288_wire_2589, c6288_wire_2588});
or_n #(2, 0, 0) OR_442 (c6288_wire_1754, {c6288_wire_689, c6288_wire_2590});
nand_n #(2, 0, 0) NAND_191 (c6288_wire_2591, {c6288_wire_67_40, c6288_wire_87_44});
notg #(0, 0) NOT_447 (c6288_wire_2592, c6288_wire_690_1);
and_n #(2, 0, 0) AND_995 (c6288_wire_2590, {c6288_wire_2592, c6288_wire_2591});
or_n #(2, 0, 0) OR_443 (c6288_wire_1759, {c6288_wire_687, c6288_wire_2593});
nand_n #(2, 0, 0) NAND_192 (c6288_wire_2594, {c6288_wire_67_41, c6288_wire_90_44});
notg #(0, 0) NOT_448 (c6288_wire_2595, c6288_wire_688_1);
and_n #(2, 0, 0) AND_996 (c6288_wire_2593, {c6288_wire_2595, c6288_wire_2594});
or_n #(2, 0, 0) OR_444 (c6288_wire_1764, {c6288_wire_685, c6288_wire_2596});
nand_n #(2, 0, 0) NAND_193 (c6288_wire_2597, {c6288_wire_67_42, c6288_wire_93_44});
notg #(0, 0) NOT_449 (c6288_wire_2598, c6288_wire_686_1);
and_n #(2, 0, 0) AND_997 (c6288_wire_2596, {c6288_wire_2598, c6288_wire_2597});
or_n #(2, 0, 0) OR_445 (c6288_wire_1769, {c6288_wire_683, c6288_wire_2599});
nand_n #(2, 0, 0) NAND_194 (c6288_wire_2600, {c6288_wire_67_43, c6288_wire_96_44});
notg #(0, 0) NOT_450 (c6288_wire_2601, c6288_wire_684_1);
and_n #(2, 0, 0) AND_998 (c6288_wire_2599, {c6288_wire_2601, c6288_wire_2600});
or_n #(2, 0, 0) OR_446 (c6288_wire_1774, {c6288_wire_681, c6288_wire_2602});
nand_n #(2, 0, 0) NAND_195 (c6288_wire_2603, {c6288_wire_67_44, c6288_wire_99_44});
notg #(0, 0) NOT_451 (c6288_wire_2604, c6288_wire_682_1);
and_n #(2, 0, 0) AND_999 (c6288_wire_2602, {c6288_wire_2604, c6288_wire_2603});
or_n #(2, 0, 0) OR_447 (c6288_wire_1711, {c6288_wire_679, c6288_wire_2605});
nand_n #(2, 0, 0) NAND_196 (c6288_wire_2606, {c6288_wire_67_45, c6288_wire_102_44});
notg #(0, 0) NOT_452 (c6288_wire_2607, c6288_wire_680_1);
and_n #(2, 0, 0) AND_1000 (c6288_wire_2605, {c6288_wire_2607, c6288_wire_2606});
or_n #(2, 0, 0) OR_448 (c6288_wire_1781, {c6288_wire_8, c6288_wire_2608});
nand_n #(2, 0, 0) NAND_197 (c6288_wire_2609, {c6288_wire_5_31, c6288_wire_6_46});
and_n #(2, 0, 0) AND_1001 (c6288_wire_2608, {c6288_wire_7, c6288_wire_2609});
or_n #(2, 0, 0) OR_449 (c6288_wire_1784, {c6288_wire_719, c6288_wire_2610});
nand_n #(2, 0, 0) NAND_198 (c6288_wire_2611, {c6288_wire_5_32, c6288_wire_105_45});
notg #(0, 0) NOT_453 (c6288_wire_2612, c6288_wire_720_1);
and_n #(2, 0, 0) AND_1002 (c6288_wire_2610, {c6288_wire_2612, c6288_wire_2611});
or_n #(2, 0, 0) OR_450 (c6288_wire_1792, {c6288_wire_717, c6288_wire_2613});
nand_n #(2, 0, 0) NAND_199 (c6288_wire_2614, {c6288_wire_5_33, c6288_wire_108_45});
notg #(0, 0) NOT_454 (c6288_wire_2615, c6288_wire_718_1);
and_n #(2, 0, 0) AND_1003 (c6288_wire_2613, {c6288_wire_2615, c6288_wire_2614});
or_n #(2, 0, 0) OR_451 (c6288_wire_1797, {c6288_wire_715, c6288_wire_2616});
nand_n #(2, 0, 0) NAND_200 (c6288_wire_2617, {c6288_wire_5_34, c6288_wire_111_45});
notg #(0, 0) NOT_455 (c6288_wire_2618, c6288_wire_716_1);
and_n #(2, 0, 0) AND_1004 (c6288_wire_2616, {c6288_wire_2618, c6288_wire_2617});
or_n #(2, 0, 0) OR_452 (c6288_wire_1802, {c6288_wire_713, c6288_wire_2619});
nand_n #(2, 0, 0) NAND_201 (c6288_wire_2620, {c6288_wire_5_35, c6288_wire_114_45});
notg #(0, 0) NOT_456 (c6288_wire_2621, c6288_wire_714_1);
and_n #(2, 0, 0) AND_1005 (c6288_wire_2619, {c6288_wire_2621, c6288_wire_2620});
or_n #(2, 0, 0) OR_453 (c6288_wire_1807, {c6288_wire_711, c6288_wire_2622});
nand_n #(2, 0, 0) NAND_202 (c6288_wire_2623, {c6288_wire_5_36, c6288_wire_117_45});
notg #(0, 0) NOT_457 (c6288_wire_2624, c6288_wire_712_1);
and_n #(2, 0, 0) AND_1006 (c6288_wire_2622, {c6288_wire_2624, c6288_wire_2623});
nor_n #(2, 0, 0) NOR_15 (c6288_wire_1968, {c6288_wire_1813_2, c6288_wire_1812_2});
or_n #(2, 0, 0) OR_454 (c6288_wire_1816, {c6288_wire_737, c6288_wire_2625});
nand_n #(2, 0, 0) NAND_203 (c6288_wire_2626, {c6288_wire_5_37, c6288_wire_78_45});
notg #(0, 0) NOT_458 (c6288_wire_2627, c6288_wire_738_1);
and_n #(2, 0, 0) AND_1007 (c6288_wire_2625, {c6288_wire_2627, c6288_wire_2626});
or_n #(2, 0, 0) OR_455 (c6288_wire_1822, {c6288_wire_735, c6288_wire_2628});
nand_n #(2, 0, 0) NAND_204 (c6288_wire_2629, {c6288_wire_5_38, c6288_wire_81_45});
notg #(0, 0) NOT_459 (c6288_wire_2630, c6288_wire_736_1);
and_n #(2, 0, 0) AND_1008 (c6288_wire_2628, {c6288_wire_2630, c6288_wire_2629});
or_n #(2, 0, 0) OR_456 (c6288_wire_1827, {c6288_wire_733, c6288_wire_2631});
nand_n #(2, 0, 0) NAND_205 (c6288_wire_2632, {c6288_wire_5_39, c6288_wire_84_45});
notg #(0, 0) NOT_460 (c6288_wire_2633, c6288_wire_734_1);
and_n #(2, 0, 0) AND_1009 (c6288_wire_2631, {c6288_wire_2633, c6288_wire_2632});
or_n #(2, 0, 0) OR_457 (c6288_wire_1832, {c6288_wire_731, c6288_wire_2634});
nand_n #(2, 0, 0) NAND_206 (c6288_wire_2635, {c6288_wire_5_40, c6288_wire_87_45});
notg #(0, 0) NOT_461 (c6288_wire_2636, c6288_wire_732_1);
and_n #(2, 0, 0) AND_1010 (c6288_wire_2634, {c6288_wire_2636, c6288_wire_2635});
or_n #(2, 0, 0) OR_458 (c6288_wire_1837, {c6288_wire_729, c6288_wire_2637});
nand_n #(2, 0, 0) NAND_207 (c6288_wire_2638, {c6288_wire_5_41, c6288_wire_90_45});
notg #(0, 0) NOT_462 (c6288_wire_2639, c6288_wire_730_1);
and_n #(2, 0, 0) AND_1011 (c6288_wire_2637, {c6288_wire_2639, c6288_wire_2638});
or_n #(2, 0, 0) OR_459 (c6288_wire_1842, {c6288_wire_727, c6288_wire_2640});
nand_n #(2, 0, 0) NAND_208 (c6288_wire_2641, {c6288_wire_5_42, c6288_wire_93_45});
notg #(0, 0) NOT_463 (c6288_wire_2642, c6288_wire_728_1);
and_n #(2, 0, 0) AND_1012 (c6288_wire_2640, {c6288_wire_2642, c6288_wire_2641});
or_n #(2, 0, 0) OR_460 (c6288_wire_1847, {c6288_wire_725, c6288_wire_2643});
nand_n #(2, 0, 0) NAND_209 (c6288_wire_2644, {c6288_wire_5_43, c6288_wire_96_45});
notg #(0, 0) NOT_464 (c6288_wire_2645, c6288_wire_726_1);
and_n #(2, 0, 0) AND_1013 (c6288_wire_2643, {c6288_wire_2645, c6288_wire_2644});
or_n #(2, 0, 0) OR_461 (c6288_wire_1852, {c6288_wire_723, c6288_wire_2646});
nand_n #(2, 0, 0) NAND_210 (c6288_wire_2647, {c6288_wire_5_44, c6288_wire_99_45});
notg #(0, 0) NOT_465 (c6288_wire_2648, c6288_wire_724_1);
and_n #(2, 0, 0) AND_1014 (c6288_wire_2646, {c6288_wire_2648, c6288_wire_2647});
or_n #(2, 0, 0) OR_462 (c6288_wire_1789, {c6288_wire_721, c6288_wire_2649});
nand_n #(2, 0, 0) NAND_211 (c6288_wire_2650, {c6288_wire_5_45, c6288_wire_102_45});
notg #(0, 0) NOT_466 (c6288_wire_2651, c6288_wire_722_1);
and_n #(2, 0, 0) AND_1015 (c6288_wire_2649, {c6288_wire_2651, c6288_wire_2650});
notg #(0, 0) NOT_467 (c6288_wire_2652, c6288_wire_833_2);
notg #(0, 0) NOT_468 (c6288_wire_2653, c6288_wire_748_2);
notg #(0, 0) NOT_469 (c6288_wire_2654, c6288_wire_757_2);
notg #(0, 0) NOT_470 (c6288_wire_2655, c6288_wire_763_2);
notg #(0, 0) NOT_471 (c6288_wire_2656, c6288_wire_769_2);
or_n #(2, 0, 0) OR_463 (c6288_wire_2015, {c6288_wire_745, c6288_wire_2657});
notg #(0, 0) NOT_472 (c6288_wire_2658, c6288_wire_2015_2);
nor_n #(2, 0, 0) NOR_16 (c6288_wire_2657, {c6288_wire_746_2, c6288_wire_31_2});
notg #(0, 0) NOT_473 (c6288_wire_2659, c6288_wire_784_2);
notg #(0, 0) NOT_474 (c6288_wire_2660, c6288_wire_791_2);
notg #(0, 0) NOT_475 (c6288_wire_2661, c6288_wire_797_2);
notg #(0, 0) NOT_476 (c6288_wire_2662, c6288_wire_803_2);
notg #(0, 0) NOT_477 (c6288_wire_2663, c6288_wire_809_2);
notg #(0, 0) NOT_478 (c6288_wire_2664, c6288_wire_815_2);
notg #(0, 0) NOT_479 (c6288_wire_2665, c6288_wire_821_2);
notg #(0, 0) NOT_480 (c6288_wire_2666, c6288_wire_827_2);
notg #(0, 0) NOT_481 (c6288_wire_2667, c6288_wire_142_2);
notg #(0, 0) NOT_482 (c6288_wire_2668, c6288_wire_140_2);
notg #(0, 0) NOT_483 (c6288_wire_2669, c6288_wire_138_2);
notg #(0, 0) NOT_484 (c6288_wire_2670, c6288_wire_136_2);
notg #(0, 0) NOT_485 (c6288_wire_2671, c6288_wire_134_2);
or_n #(2, 0, 0) OR_464 (c6288_wire_160, {c6288_wire_836, c6288_wire_2672});
notg #(0, 0) NOT_486 (c6288_wire_2673, c6288_wire_160_2);
nor_n #(2, 0, 0) NOR_17 (c6288_wire_2672, {c6288_wire_837_2, c6288_wire_11_2});
notg #(0, 0) NOT_487 (c6288_wire_2674, c6288_wire_158_2);
notg #(0, 0) NOT_488 (c6288_wire_2675, c6288_wire_156_2);
notg #(0, 0) NOT_489 (c6288_wire_2676, c6288_wire_154_2);
notg #(0, 0) NOT_490 (c6288_wire_2677, c6288_wire_152_2);
notg #(0, 0) NOT_491 (c6288_wire_2678, c6288_wire_150_2);
notg #(0, 0) NOT_492 (c6288_wire_2679, c6288_wire_148_2);
notg #(0, 0) NOT_493 (c6288_wire_2680, c6288_wire_146_2);
notg #(0, 0) NOT_494 (c6288_wire_2681, c6288_wire_144_2);
notg #(0, 0) NOT_495 (c6288_wire_2682, c6288_wire_184_2);
notg #(0, 0) NOT_496 (c6288_wire_2683, c6288_wire_182_2);
notg #(0, 0) NOT_497 (c6288_wire_2684, c6288_wire_180_2);
notg #(0, 0) NOT_498 (c6288_wire_2685, c6288_wire_178_2);
notg #(0, 0) NOT_499 (c6288_wire_2686, c6288_wire_176_2);
or_n #(2, 0, 0) OR_465 (c6288_wire_202, {c6288_wire_917, c6288_wire_2687});
notg #(0, 0) NOT_500 (c6288_wire_2688, c6288_wire_202_2);
nor_n #(2, 0, 0) NOR_18 (c6288_wire_2687, {c6288_wire_918_2, c6288_wire_16_2});
notg #(0, 0) NOT_501 (c6288_wire_2689, c6288_wire_200_2);
notg #(0, 0) NOT_502 (c6288_wire_2690, c6288_wire_198_2);
notg #(0, 0) NOT_503 (c6288_wire_2691, c6288_wire_196_2);
notg #(0, 0) NOT_504 (c6288_wire_2692, c6288_wire_194_2);
notg #(0, 0) NOT_505 (c6288_wire_2693, c6288_wire_192_2);
notg #(0, 0) NOT_506 (c6288_wire_2694, c6288_wire_190_2);
notg #(0, 0) NOT_507 (c6288_wire_2695, c6288_wire_188_2);
notg #(0, 0) NOT_508 (c6288_wire_2696, c6288_wire_186_2);
notg #(0, 0) NOT_509 (c6288_wire_2697, c6288_wire_226_2);
notg #(0, 0) NOT_510 (c6288_wire_2698, c6288_wire_224_2);
notg #(0, 0) NOT_511 (c6288_wire_2699, c6288_wire_222_2);
notg #(0, 0) NOT_512 (c6288_wire_2700, c6288_wire_220_2);
notg #(0, 0) NOT_513 (c6288_wire_2701, c6288_wire_218_2);
or_n #(2, 0, 0) OR_466 (c6288_wire_244, {c6288_wire_995, c6288_wire_2702});
notg #(0, 0) NOT_514 (c6288_wire_2703, c6288_wire_244_2);
nor_n #(2, 0, 0) NOR_19 (c6288_wire_2702, {c6288_wire_996_2, c6288_wire_21_2});
notg #(0, 0) NOT_515 (c6288_wire_2704, c6288_wire_242_2);
notg #(0, 0) NOT_516 (c6288_wire_2705, c6288_wire_240_2);
notg #(0, 0) NOT_517 (c6288_wire_2706, c6288_wire_238_2);
notg #(0, 0) NOT_518 (c6288_wire_2707, c6288_wire_236_2);
notg #(0, 0) NOT_519 (c6288_wire_2708, c6288_wire_234_2);
notg #(0, 0) NOT_520 (c6288_wire_2709, c6288_wire_232_2);
notg #(0, 0) NOT_521 (c6288_wire_2710, c6288_wire_230_2);
notg #(0, 0) NOT_522 (c6288_wire_2711, c6288_wire_228_2);
notg #(0, 0) NOT_523 (c6288_wire_2712, c6288_wire_268_2);
notg #(0, 0) NOT_524 (c6288_wire_2713, c6288_wire_266_2);
notg #(0, 0) NOT_525 (c6288_wire_2714, c6288_wire_264_2);
notg #(0, 0) NOT_526 (c6288_wire_2715, c6288_wire_262_2);
notg #(0, 0) NOT_527 (c6288_wire_2716, c6288_wire_260_2);
notg #(0, 0) NOT_528 (c6288_wire_2717, c6288_wire_286_2);
or_n #(2, 0, 0) OR_467 (c6288_wire_284, {c6288_wire_1107, c6288_wire_2718});
notg #(0, 0) NOT_529 (c6288_wire_2719, c6288_wire_284_2);
nor_n #(2, 0, 0) NOR_20 (c6288_wire_2718, {c6288_wire_1109_2, c6288_wire_1108_2});
notg #(0, 0) NOT_530 (c6288_wire_2720, c6288_wire_282_2);
notg #(0, 0) NOT_531 (c6288_wire_2721, c6288_wire_280_2);
notg #(0, 0) NOT_532 (c6288_wire_2722, c6288_wire_278_2);
notg #(0, 0) NOT_533 (c6288_wire_2723, c6288_wire_276_2);
notg #(0, 0) NOT_534 (c6288_wire_2724, c6288_wire_274_2);
notg #(0, 0) NOT_535 (c6288_wire_2725, c6288_wire_272_2);
notg #(0, 0) NOT_536 (c6288_wire_2726, c6288_wire_270_2);
notg #(0, 0) NOT_537 (c6288_wire_2727, c6288_wire_311_2);
or_n #(2, 0, 0) OR_468 (c6288_wire_311, {c6288_wire_2728, c6288_wire_1231});
nand_n #(2, 0, 0) NAND_212 (c6288_wire_1232, {c6288_wire_330_31, c6288_wire_102_46});
and_n #(2, 0, 0) AND_1016 (c6288_wire_2728, {c6288_wire_347, c6288_wire_1230});
notg #(0, 0) NOT_538 (c6288_wire_2729, c6288_wire_309_2);
or_n #(2, 0, 0) OR_469 (c6288_wire_309, {c6288_wire_2730, c6288_wire_1157});
nand_n #(2, 0, 0) NAND_213 (c6288_wire_1158, {c6288_wire_330_32, c6288_wire_105_46});
and_n #(2, 0, 0) AND_1017 (c6288_wire_2730, {c6288_wire_346, c6288_wire_1156});
notg #(0, 0) NOT_539 (c6288_wire_2731, c6288_wire_307_2);
or_n #(2, 0, 0) OR_470 (c6288_wire_307, {c6288_wire_2732, c6288_wire_1163});
nand_n #(2, 0, 0) NAND_214 (c6288_wire_1164, {c6288_wire_330_33, c6288_wire_108_46});
and_n #(2, 0, 0) AND_1018 (c6288_wire_2732, {c6288_wire_345, c6288_wire_1162});
notg #(0, 0) NOT_540 (c6288_wire_2733, c6288_wire_305_2);
or_n #(2, 0, 0) OR_471 (c6288_wire_305, {c6288_wire_2734, c6288_wire_1169});
nand_n #(2, 0, 0) NAND_215 (c6288_wire_1170, {c6288_wire_330_34, c6288_wire_111_46});
and_n #(2, 0, 0) AND_1019 (c6288_wire_2734, {c6288_wire_344, c6288_wire_1168});
notg #(0, 0) NOT_541 (c6288_wire_2735, c6288_wire_303_2);
or_n #(2, 0, 0) OR_472 (c6288_wire_303, {c6288_wire_2736, c6288_wire_1175});
nand_n #(2, 0, 0) NAND_216 (c6288_wire_1176, {c6288_wire_330_35, c6288_wire_114_46});
and_n #(2, 0, 0) AND_1020 (c6288_wire_2736, {c6288_wire_343, c6288_wire_1174});
or_n #(2, 0, 0) OR_473 (c6288_wire_1104, {c6288_wire_2737, c6288_wire_1180});
nand_n #(2, 0, 0) NAND_217 (c6288_wire_1181, {c6288_wire_330_36, c6288_wire_117_46});
and_n #(2, 0, 0) AND_1021 (c6288_wire_2737, {c6288_wire_342, c6288_wire_1179});
notg #(0, 0) NOT_542 (c6288_wire_2738, c6288_wire_2230_2);
and_n #(2, 0, 0) AND_1022 (c6288_wire_2230, {c6288_wire_355, c6288_wire_2739});
nand_n #(2, 0, 0) NAND_218 (c6288_wire_2739, {c6288_wire_25_44, c6288_wire_3_17});
notg #(0, 0) NOT_543 (c6288_wire_2740, c6288_wire_327_2);
nand_n #(2, 0, 0) NAND_219 (c6288_wire_744, {c6288_wire_6_47, c6288_wire_740_3});
and_n #(2, 0, 0) AND_1023 (c6288_wire_2741, {c6288_wire_741, c6288_wire_742});
or_n #(2, 0, 0) OR_474 (c6288_wire_360, {c6288_wire_2741, c6288_wire_743});
notg #(0, 0) NOT_544 (c6288_wire_2742, c6288_wire_325_2);
or_n #(2, 0, 0) OR_475 (c6288_wire_325, {c6288_wire_2743, c6288_wire_1190});
nand_n #(2, 0, 0) NAND_220 (c6288_wire_1191, {c6288_wire_330_37, c6288_wire_81_46});
and_n #(2, 0, 0) AND_1024 (c6288_wire_2743, {c6288_wire_354, c6288_wire_1189});
notg #(0, 0) NOT_545 (c6288_wire_2744, c6288_wire_323_2);
or_n #(2, 0, 0) OR_476 (c6288_wire_323, {c6288_wire_2745, c6288_wire_1196});
nand_n #(2, 0, 0) NAND_221 (c6288_wire_1197, {c6288_wire_330_38, c6288_wire_84_46});
and_n #(2, 0, 0) AND_1025 (c6288_wire_2745, {c6288_wire_353, c6288_wire_1195});
notg #(0, 0) NOT_546 (c6288_wire_2746, c6288_wire_321_2);
or_n #(2, 0, 0) OR_477 (c6288_wire_321, {c6288_wire_2747, c6288_wire_1202});
nand_n #(2, 0, 0) NAND_222 (c6288_wire_1203, {c6288_wire_330_39, c6288_wire_87_46});
and_n #(2, 0, 0) AND_1026 (c6288_wire_2747, {c6288_wire_352, c6288_wire_1201});
notg #(0, 0) NOT_547 (c6288_wire_2748, c6288_wire_319_2);
or_n #(2, 0, 0) OR_478 (c6288_wire_319, {c6288_wire_2749, c6288_wire_1208});
nand_n #(2, 0, 0) NAND_223 (c6288_wire_1209, {c6288_wire_330_40, c6288_wire_90_46});
and_n #(2, 0, 0) AND_1027 (c6288_wire_2749, {c6288_wire_351, c6288_wire_1207});
notg #(0, 0) NOT_548 (c6288_wire_2750, c6288_wire_317_2);
or_n #(2, 0, 0) OR_479 (c6288_wire_317, {c6288_wire_2751, c6288_wire_1214});
nand_n #(2, 0, 0) NAND_224 (c6288_wire_1215, {c6288_wire_330_41, c6288_wire_93_46});
and_n #(2, 0, 0) AND_1028 (c6288_wire_2751, {c6288_wire_350, c6288_wire_1213});
notg #(0, 0) NOT_549 (c6288_wire_2752, c6288_wire_315_2);
or_n #(2, 0, 0) OR_480 (c6288_wire_315, {c6288_wire_2753, c6288_wire_1220});
nand_n #(2, 0, 0) NAND_225 (c6288_wire_1221, {c6288_wire_330_42, c6288_wire_96_46});
and_n #(2, 0, 0) AND_1029 (c6288_wire_2753, {c6288_wire_349, c6288_wire_1219});
notg #(0, 0) NOT_550 (c6288_wire_2754, c6288_wire_313_2);
or_n #(2, 0, 0) OR_481 (c6288_wire_313, {c6288_wire_2755, c6288_wire_1226});
nand_n #(2, 0, 0) NAND_226 (c6288_wire_1227, {c6288_wire_330_43, c6288_wire_99_46});
and_n #(2, 0, 0) AND_1030 (c6288_wire_2755, {c6288_wire_348, c6288_wire_1225});
notg #(0, 0) NOT_551 (c6288_wire_2756, c6288_wire_384_2);
notg #(0, 0) NOT_552 (c6288_wire_2757, c6288_wire_382_2);
notg #(0, 0) NOT_553 (c6288_wire_2758, c6288_wire_380_2);
notg #(0, 0) NOT_554 (c6288_wire_2759, c6288_wire_378_2);
notg #(0, 0) NOT_555 (c6288_wire_2760, c6288_wire_376_2);
or_n #(2, 0, 0) OR_482 (c6288_wire_402, {c6288_wire_1233, c6288_wire_2761});
notg #(0, 0) NOT_556 (c6288_wire_2762, c6288_wire_402_2);
nor_n #(2, 0, 0) NOR_21 (c6288_wire_2761, {c6288_wire_1234_2, c6288_wire_38_2});
notg #(0, 0) NOT_557 (c6288_wire_2763, c6288_wire_400_2);
notg #(0, 0) NOT_558 (c6288_wire_2764, c6288_wire_398_2);
notg #(0, 0) NOT_559 (c6288_wire_2765, c6288_wire_396_2);
notg #(0, 0) NOT_560 (c6288_wire_2766, c6288_wire_394_2);
notg #(0, 0) NOT_561 (c6288_wire_2767, c6288_wire_392_2);
notg #(0, 0) NOT_562 (c6288_wire_2768, c6288_wire_390_2);
notg #(0, 0) NOT_563 (c6288_wire_2769, c6288_wire_388_2);
notg #(0, 0) NOT_564 (c6288_wire_2770, c6288_wire_386_2);
notg #(0, 0) NOT_565 (c6288_wire_2771, c6288_wire_426_2);
notg #(0, 0) NOT_566 (c6288_wire_2772, c6288_wire_424_2);
notg #(0, 0) NOT_567 (c6288_wire_2773, c6288_wire_422_2);
notg #(0, 0) NOT_568 (c6288_wire_2774, c6288_wire_420_2);
notg #(0, 0) NOT_569 (c6288_wire_2775, c6288_wire_418_2);
or_n #(2, 0, 0) OR_483 (c6288_wire_444, {c6288_wire_1312, c6288_wire_2776});
notg #(0, 0) NOT_570 (c6288_wire_2777, c6288_wire_444_2);
nor_n #(2, 0, 0) NOR_22 (c6288_wire_2776, {c6288_wire_1313_2, c6288_wire_43_2});
notg #(0, 0) NOT_571 (c6288_wire_2778, c6288_wire_442_2);
notg #(0, 0) NOT_572 (c6288_wire_2779, c6288_wire_440_2);
notg #(0, 0) NOT_573 (c6288_wire_2780, c6288_wire_438_2);
notg #(0, 0) NOT_574 (c6288_wire_2781, c6288_wire_436_2);
notg #(0, 0) NOT_575 (c6288_wire_2782, c6288_wire_434_2);
notg #(0, 0) NOT_576 (c6288_wire_2783, c6288_wire_432_2);
notg #(0, 0) NOT_577 (c6288_wire_2784, c6288_wire_430_2);
notg #(0, 0) NOT_578 (c6288_wire_2785, c6288_wire_428_2);
notg #(0, 0) NOT_579 (c6288_wire_2786, c6288_wire_468_2);
notg #(0, 0) NOT_580 (c6288_wire_2787, c6288_wire_466_2);
notg #(0, 0) NOT_581 (c6288_wire_2788, c6288_wire_464_2);
notg #(0, 0) NOT_582 (c6288_wire_2789, c6288_wire_462_2);
notg #(0, 0) NOT_583 (c6288_wire_2790, c6288_wire_460_2);
or_n #(2, 0, 0) OR_484 (c6288_wire_486, {c6288_wire_1390, c6288_wire_2791});
notg #(0, 0) NOT_584 (c6288_wire_2792, c6288_wire_486_2);
nor_n #(2, 0, 0) NOR_23 (c6288_wire_2791, {c6288_wire_1391_2, c6288_wire_48_2});
notg #(0, 0) NOT_585 (c6288_wire_2793, c6288_wire_484_2);
notg #(0, 0) NOT_586 (c6288_wire_2794, c6288_wire_482_2);
notg #(0, 0) NOT_587 (c6288_wire_2795, c6288_wire_480_2);
notg #(0, 0) NOT_588 (c6288_wire_2796, c6288_wire_478_2);
notg #(0, 0) NOT_589 (c6288_wire_2797, c6288_wire_476_2);
notg #(0, 0) NOT_590 (c6288_wire_2798, c6288_wire_474_2);
notg #(0, 0) NOT_591 (c6288_wire_2799, c6288_wire_472_2);
notg #(0, 0) NOT_592 (c6288_wire_2800, c6288_wire_470_2);
notg #(0, 0) NOT_593 (c6288_wire_2801, c6288_wire_510_2);
notg #(0, 0) NOT_594 (c6288_wire_2802, c6288_wire_508_2);
notg #(0, 0) NOT_595 (c6288_wire_2803, c6288_wire_506_2);
notg #(0, 0) NOT_596 (c6288_wire_2804, c6288_wire_504_2);
notg #(0, 0) NOT_597 (c6288_wire_2805, c6288_wire_502_2);
or_n #(2, 0, 0) OR_485 (c6288_wire_528, {c6288_wire_1468, c6288_wire_2806});
notg #(0, 0) NOT_598 (c6288_wire_2807, c6288_wire_528_2);
nor_n #(2, 0, 0) NOR_24 (c6288_wire_2806, {c6288_wire_1469_2, c6288_wire_53_2});
notg #(0, 0) NOT_599 (c6288_wire_2808, c6288_wire_526_2);
notg #(0, 0) NOT_600 (c6288_wire_2809, c6288_wire_524_2);
notg #(0, 0) NOT_601 (c6288_wire_2810, c6288_wire_522_2);
notg #(0, 0) NOT_602 (c6288_wire_2811, c6288_wire_520_2);
notg #(0, 0) NOT_603 (c6288_wire_2812, c6288_wire_518_2);
notg #(0, 0) NOT_604 (c6288_wire_2813, c6288_wire_516_2);
notg #(0, 0) NOT_605 (c6288_wire_2814, c6288_wire_514_2);
notg #(0, 0) NOT_606 (c6288_wire_2815, c6288_wire_512_2);
notg #(0, 0) NOT_607 (c6288_wire_2816, c6288_wire_552_2);
notg #(0, 0) NOT_608 (c6288_wire_2817, c6288_wire_550_2);
notg #(0, 0) NOT_609 (c6288_wire_2818, c6288_wire_548_2);
notg #(0, 0) NOT_610 (c6288_wire_2819, c6288_wire_546_2);
notg #(0, 0) NOT_611 (c6288_wire_2820, c6288_wire_544_2);
or_n #(2, 0, 0) OR_486 (c6288_wire_570, {c6288_wire_1546, c6288_wire_2821});
notg #(0, 0) NOT_612 (c6288_wire_2822, c6288_wire_570_2);
nor_n #(2, 0, 0) NOR_25 (c6288_wire_2821, {c6288_wire_1547_2, c6288_wire_58_2});
notg #(0, 0) NOT_613 (c6288_wire_2823, c6288_wire_568_2);
notg #(0, 0) NOT_614 (c6288_wire_2824, c6288_wire_566_2);
notg #(0, 0) NOT_615 (c6288_wire_2825, c6288_wire_564_2);
notg #(0, 0) NOT_616 (c6288_wire_2826, c6288_wire_562_2);
notg #(0, 0) NOT_617 (c6288_wire_2827, c6288_wire_560_2);
notg #(0, 0) NOT_618 (c6288_wire_2828, c6288_wire_558_2);
notg #(0, 0) NOT_619 (c6288_wire_2829, c6288_wire_556_2);
notg #(0, 0) NOT_620 (c6288_wire_2830, c6288_wire_554_2);
notg #(0, 0) NOT_621 (c6288_wire_2831, c6288_wire_594_2);
notg #(0, 0) NOT_622 (c6288_wire_2832, c6288_wire_592_2);
notg #(0, 0) NOT_623 (c6288_wire_2833, c6288_wire_590_2);
notg #(0, 0) NOT_624 (c6288_wire_2834, c6288_wire_588_2);
notg #(0, 0) NOT_625 (c6288_wire_2835, c6288_wire_586_2);
or_n #(2, 0, 0) OR_487 (c6288_wire_612, {c6288_wire_1624, c6288_wire_2836});
notg #(0, 0) NOT_626 (c6288_wire_2837, c6288_wire_612_2);
nor_n #(2, 0, 0) NOR_26 (c6288_wire_2836, {c6288_wire_1625_2, c6288_wire_63_2});
notg #(0, 0) NOT_627 (c6288_wire_2838, c6288_wire_610_2);
notg #(0, 0) NOT_628 (c6288_wire_2839, c6288_wire_608_2);
notg #(0, 0) NOT_629 (c6288_wire_2840, c6288_wire_606_2);
notg #(0, 0) NOT_630 (c6288_wire_2841, c6288_wire_604_2);
notg #(0, 0) NOT_631 (c6288_wire_2842, c6288_wire_602_2);
notg #(0, 0) NOT_632 (c6288_wire_2843, c6288_wire_600_2);
notg #(0, 0) NOT_633 (c6288_wire_2844, c6288_wire_598_2);
notg #(0, 0) NOT_634 (c6288_wire_2845, c6288_wire_596_2);
notg #(0, 0) NOT_635 (c6288_wire_2846, c6288_wire_636_2);
notg #(0, 0) NOT_636 (c6288_wire_2847, c6288_wire_634_2);
notg #(0, 0) NOT_637 (c6288_wire_2848, c6288_wire_632_2);
notg #(0, 0) NOT_638 (c6288_wire_2849, c6288_wire_630_2);
notg #(0, 0) NOT_639 (c6288_wire_2850, c6288_wire_628_2);
or_n #(2, 0, 0) OR_488 (c6288_wire_654, {c6288_wire_1702, c6288_wire_2851});
notg #(0, 0) NOT_640 (c6288_wire_2852, c6288_wire_654_2);
nor_n #(2, 0, 0) NOR_27 (c6288_wire_2851, {c6288_wire_1703_2, c6288_wire_68_2});
notg #(0, 0) NOT_641 (c6288_wire_2853, c6288_wire_652_2);
notg #(0, 0) NOT_642 (c6288_wire_2854, c6288_wire_650_2);
notg #(0, 0) NOT_643 (c6288_wire_2855, c6288_wire_648_2);
notg #(0, 0) NOT_644 (c6288_wire_2856, c6288_wire_646_2);
notg #(0, 0) NOT_645 (c6288_wire_2857, c6288_wire_644_2);
notg #(0, 0) NOT_646 (c6288_wire_2858, c6288_wire_642_2);
notg #(0, 0) NOT_647 (c6288_wire_2859, c6288_wire_640_2);
notg #(0, 0) NOT_648 (c6288_wire_2860, c6288_wire_638_2);
notg #(0, 0) NOT_649 (c6288_wire_2861, c6288_wire_678_2);
notg #(0, 0) NOT_650 (c6288_wire_2862, c6288_wire_676_2);
notg #(0, 0) NOT_651 (c6288_wire_2863, c6288_wire_674_2);
notg #(0, 0) NOT_652 (c6288_wire_2864, c6288_wire_672_2);
notg #(0, 0) NOT_653 (c6288_wire_2865, c6288_wire_670_2);
or_n #(2, 0, 0) OR_489 (c6288_wire_696, {c6288_wire_1780, c6288_wire_2866});
notg #(0, 0) NOT_654 (c6288_wire_2867, c6288_wire_696_2);
nor_n #(2, 0, 0) NOR_28 (c6288_wire_2866, {c6288_wire_1781_2, c6288_wire_72_2});
notg #(0, 0) NOT_655 (c6288_wire_2868, c6288_wire_694_2);
notg #(0, 0) NOT_656 (c6288_wire_2869, c6288_wire_692_2);
notg #(0, 0) NOT_657 (c6288_wire_2870, c6288_wire_690_2);
notg #(0, 0) NOT_658 (c6288_wire_2871, c6288_wire_688_2);
notg #(0, 0) NOT_659 (c6288_wire_2872, c6288_wire_686_2);
notg #(0, 0) NOT_660 (c6288_wire_2873, c6288_wire_684_2);
notg #(0, 0) NOT_661 (c6288_wire_2874, c6288_wire_682_2);
notg #(0, 0) NOT_662 (c6288_wire_2875, c6288_wire_680_2);
notg #(0, 0) NOT_663 (c6288_wire_2876, c6288_wire_720_2);
notg #(0, 0) NOT_664 (c6288_wire_2877, c6288_wire_718_2);
notg #(0, 0) NOT_665 (c6288_wire_2878, c6288_wire_716_2);
notg #(0, 0) NOT_666 (c6288_wire_2879, c6288_wire_714_2);
notg #(0, 0) NOT_667 (c6288_wire_2880, c6288_wire_712_2);
or_n #(2, 0, 0) OR_490 (c6288_wire_738, {c6288_wire_1858, c6288_wire_2881});
notg #(0, 0) NOT_668 (c6288_wire_2882, c6288_wire_738_2);
nor_n #(2, 0, 0) NOR_29 (c6288_wire_2881, {c6288_wire_1859_2, c6288_wire_4_2});
notg #(0, 0) NOT_669 (c6288_wire_2883, c6288_wire_736_2);
notg #(0, 0) NOT_670 (c6288_wire_2884, c6288_wire_734_2);
notg #(0, 0) NOT_671 (c6288_wire_2885, c6288_wire_732_2);
notg #(0, 0) NOT_672 (c6288_wire_2886, c6288_wire_730_2);
notg #(0, 0) NOT_673 (c6288_wire_2887, c6288_wire_728_2);
notg #(0, 0) NOT_674 (c6288_wire_2888, c6288_wire_726_2);
notg #(0, 0) NOT_675 (c6288_wire_2889, c6288_wire_724_2);
notg #(0, 0) NOT_676 (c6288_wire_2890, c6288_wire_722_2);
or_n #(2, 0, 0) OR_491 (c6288_wire_756, {c6288_wire_104, c6288_wire_2652});
or_n #(2, 0, 0) OR_492 (c6288_wire_762, {c6288_wire_107, c6288_wire_2653});
or_n #(2, 0, 0) OR_493 (c6288_wire_768, {c6288_wire_110, c6288_wire_2654});
or_n #(2, 0, 0) OR_494 (c6288_wire_774, {c6288_wire_113, c6288_wire_2655});
or_n #(2, 0, 0) OR_495 (c6288_wire_779, {c6288_wire_116, c6288_wire_2656});
or_n #(2, 0, 0) OR_496 (c6288_wire_790, {c6288_wire_77, c6288_wire_2658});
or_n #(2, 0, 0) OR_497 (c6288_wire_796, {c6288_wire_80, c6288_wire_2659});
or_n #(2, 0, 0) OR_498 (c6288_wire_802, {c6288_wire_83, c6288_wire_2660});
or_n #(2, 0, 0) OR_499 (c6288_wire_808, {c6288_wire_86, c6288_wire_2661});
or_n #(2, 0, 0) OR_500 (c6288_wire_814, {c6288_wire_89, c6288_wire_2662});
or_n #(2, 0, 0) OR_501 (c6288_wire_820, {c6288_wire_92, c6288_wire_2663});
or_n #(2, 0, 0) OR_502 (c6288_wire_826, {c6288_wire_95, c6288_wire_2664});
or_n #(2, 0, 0) OR_503 (c6288_wire_832, {c6288_wire_98, c6288_wire_2665});
or_n #(2, 0, 0) OR_504 (c6288_wire_835, {c6288_wire_101, c6288_wire_2666});
or_n #(2, 0, 0) OR_505 (c6288_wire_846, {c6288_wire_128, c6288_wire_2667});
or_n #(2, 0, 0) OR_506 (c6288_wire_851, {c6288_wire_129, c6288_wire_2668});
or_n #(2, 0, 0) OR_507 (c6288_wire_856, {c6288_wire_130, c6288_wire_2669});
or_n #(2, 0, 0) OR_508 (c6288_wire_861, {c6288_wire_131, c6288_wire_2670});
or_n #(2, 0, 0) OR_509 (c6288_wire_867, {c6288_wire_132, c6288_wire_2671});
or_n #(2, 0, 0) OR_510 (c6288_wire_879, {c6288_wire_119, c6288_wire_2673});
or_n #(2, 0, 0) OR_511 (c6288_wire_884, {c6288_wire_120, c6288_wire_2674});
or_n #(2, 0, 0) OR_512 (c6288_wire_889, {c6288_wire_121, c6288_wire_2675});
or_n #(2, 0, 0) OR_513 (c6288_wire_894, {c6288_wire_122, c6288_wire_2676});
or_n #(2, 0, 0) OR_514 (c6288_wire_899, {c6288_wire_123, c6288_wire_2677});
or_n #(2, 0, 0) OR_515 (c6288_wire_904, {c6288_wire_124, c6288_wire_2678});
or_n #(2, 0, 0) OR_516 (c6288_wire_909, {c6288_wire_125, c6288_wire_2679});
or_n #(2, 0, 0) OR_517 (c6288_wire_914, {c6288_wire_126, c6288_wire_2680});
or_n #(2, 0, 0) OR_518 (c6288_wire_916, {c6288_wire_127, c6288_wire_2681});
or_n #(2, 0, 0) OR_519 (c6288_wire_927, {c6288_wire_170, c6288_wire_2682});
or_n #(2, 0, 0) OR_520 (c6288_wire_932, {c6288_wire_171, c6288_wire_2683});
or_n #(2, 0, 0) OR_521 (c6288_wire_937, {c6288_wire_172, c6288_wire_2684});
or_n #(2, 0, 0) OR_522 (c6288_wire_942, {c6288_wire_173, c6288_wire_2685});
or_n #(2, 0, 0) OR_523 (c6288_wire_947, {c6288_wire_174, c6288_wire_2686});
or_n #(2, 0, 0) OR_524 (c6288_wire_957, {c6288_wire_161, c6288_wire_2688});
or_n #(2, 0, 0) OR_525 (c6288_wire_962, {c6288_wire_162, c6288_wire_2689});
or_n #(2, 0, 0) OR_526 (c6288_wire_967, {c6288_wire_163, c6288_wire_2690});
or_n #(2, 0, 0) OR_527 (c6288_wire_972, {c6288_wire_164, c6288_wire_2691});
or_n #(2, 0, 0) OR_528 (c6288_wire_977, {c6288_wire_165, c6288_wire_2692});
or_n #(2, 0, 0) OR_529 (c6288_wire_982, {c6288_wire_166, c6288_wire_2693});
or_n #(2, 0, 0) OR_530 (c6288_wire_987, {c6288_wire_167, c6288_wire_2694});
or_n #(2, 0, 0) OR_531 (c6288_wire_992, {c6288_wire_168, c6288_wire_2695});
or_n #(2, 0, 0) OR_532 (c6288_wire_994, {c6288_wire_169, c6288_wire_2696});
or_n #(2, 0, 0) OR_533 (c6288_wire_1005, {c6288_wire_212, c6288_wire_2697});
or_n #(2, 0, 0) OR_534 (c6288_wire_1010, {c6288_wire_213, c6288_wire_2698});
or_n #(2, 0, 0) OR_535 (c6288_wire_1015, {c6288_wire_214, c6288_wire_2699});
or_n #(2, 0, 0) OR_536 (c6288_wire_1020, {c6288_wire_215, c6288_wire_2700});
or_n #(2, 0, 0) OR_537 (c6288_wire_1025, {c6288_wire_216, c6288_wire_2701});
or_n #(2, 0, 0) OR_538 (c6288_wire_1035, {c6288_wire_203, c6288_wire_2703});
or_n #(2, 0, 0) OR_539 (c6288_wire_1040, {c6288_wire_204, c6288_wire_2704});
or_n #(2, 0, 0) OR_540 (c6288_wire_1045, {c6288_wire_205, c6288_wire_2705});
or_n #(2, 0, 0) OR_541 (c6288_wire_1050, {c6288_wire_206, c6288_wire_2706});
or_n #(2, 0, 0) OR_542 (c6288_wire_1055, {c6288_wire_207, c6288_wire_2707});
or_n #(2, 0, 0) OR_543 (c6288_wire_1060, {c6288_wire_208, c6288_wire_2708});
or_n #(2, 0, 0) OR_544 (c6288_wire_1065, {c6288_wire_209, c6288_wire_2709});
or_n #(2, 0, 0) OR_545 (c6288_wire_1070, {c6288_wire_210, c6288_wire_2710});
or_n #(2, 0, 0) OR_546 (c6288_wire_1072, {c6288_wire_211, c6288_wire_2711});
or_n #(2, 0, 0) OR_547 (c6288_wire_1081, {c6288_wire_254, c6288_wire_2712});
or_n #(2, 0, 0) OR_548 (c6288_wire_1086, {c6288_wire_255, c6288_wire_2713});
or_n #(2, 0, 0) OR_549 (c6288_wire_1091, {c6288_wire_256, c6288_wire_2714});
or_n #(2, 0, 0) OR_550 (c6288_wire_1096, {c6288_wire_257, c6288_wire_2715});
or_n #(2, 0, 0) OR_551 (c6288_wire_1101, {c6288_wire_258, c6288_wire_2716});
or_n #(2, 0, 0) OR_552 (c6288_wire_1114, {c6288_wire_245, c6288_wire_2717});
or_n #(2, 0, 0) OR_553 (c6288_wire_1119, {c6288_wire_246, c6288_wire_2719});
or_n #(2, 0, 0) OR_554 (c6288_wire_1124, {c6288_wire_247, c6288_wire_2720});
or_n #(2, 0, 0) OR_555 (c6288_wire_1129, {c6288_wire_248, c6288_wire_2721});
or_n #(2, 0, 0) OR_556 (c6288_wire_1134, {c6288_wire_249, c6288_wire_2722});
or_n #(2, 0, 0) OR_557 (c6288_wire_1139, {c6288_wire_250, c6288_wire_2723});
or_n #(2, 0, 0) OR_558 (c6288_wire_1144, {c6288_wire_251, c6288_wire_2724});
or_n #(2, 0, 0) OR_559 (c6288_wire_1149, {c6288_wire_252, c6288_wire_2725});
or_n #(2, 0, 0) OR_560 (c6288_wire_1151, {c6288_wire_253, c6288_wire_2726});
or_n #(2, 0, 0) OR_561 (c6288_wire_1154, {c6288_wire_297, c6288_wire_2727});
or_n #(2, 0, 0) OR_562 (c6288_wire_1160, {c6288_wire_298, c6288_wire_2729});
or_n #(2, 0, 0) OR_563 (c6288_wire_1166, {c6288_wire_299, c6288_wire_2731});
or_n #(2, 0, 0) OR_564 (c6288_wire_1172, {c6288_wire_300, c6288_wire_2733});
or_n #(2, 0, 0) OR_565 (c6288_wire_1178, {c6288_wire_301, c6288_wire_2735});
or_n #(2, 0, 0) OR_566 (c6288_wire_740, {c6288_wire_287, c6288_wire_2738});
or_n #(2, 0, 0) OR_567 (c6288_wire_1187, {c6288_wire_289, c6288_wire_2740});
or_n #(2, 0, 0) OR_568 (c6288_wire_1193, {c6288_wire_290, c6288_wire_2742});
or_n #(2, 0, 0) OR_569 (c6288_wire_1199, {c6288_wire_291, c6288_wire_2744});
or_n #(2, 0, 0) OR_570 (c6288_wire_1205, {c6288_wire_292, c6288_wire_2746});
or_n #(2, 0, 0) OR_571 (c6288_wire_1211, {c6288_wire_293, c6288_wire_2748});
or_n #(2, 0, 0) OR_572 (c6288_wire_1217, {c6288_wire_294, c6288_wire_2750});
or_n #(2, 0, 0) OR_573 (c6288_wire_1223, {c6288_wire_295, c6288_wire_2752});
or_n #(2, 0, 0) OR_574 (c6288_wire_1229, {c6288_wire_296, c6288_wire_2754});
or_n #(2, 0, 0) OR_575 (c6288_wire_1243, {c6288_wire_370, c6288_wire_2756});
or_n #(2, 0, 0) OR_576 (c6288_wire_1248, {c6288_wire_371, c6288_wire_2757});
or_n #(2, 0, 0) OR_577 (c6288_wire_1253, {c6288_wire_372, c6288_wire_2758});
or_n #(2, 0, 0) OR_578 (c6288_wire_1258, {c6288_wire_373, c6288_wire_2759});
or_n #(2, 0, 0) OR_579 (c6288_wire_1263, {c6288_wire_374, c6288_wire_2760});
or_n #(2, 0, 0) OR_580 (c6288_wire_1274, {c6288_wire_361, c6288_wire_2762});
or_n #(2, 0, 0) OR_581 (c6288_wire_1279, {c6288_wire_362, c6288_wire_2763});
or_n #(2, 0, 0) OR_582 (c6288_wire_1284, {c6288_wire_363, c6288_wire_2764});
or_n #(2, 0, 0) OR_583 (c6288_wire_1289, {c6288_wire_364, c6288_wire_2765});
or_n #(2, 0, 0) OR_584 (c6288_wire_1294, {c6288_wire_365, c6288_wire_2766});
or_n #(2, 0, 0) OR_585 (c6288_wire_1299, {c6288_wire_366, c6288_wire_2767});
or_n #(2, 0, 0) OR_586 (c6288_wire_1304, {c6288_wire_367, c6288_wire_2768});
or_n #(2, 0, 0) OR_587 (c6288_wire_1309, {c6288_wire_368, c6288_wire_2769});
or_n #(2, 0, 0) OR_588 (c6288_wire_1311, {c6288_wire_369, c6288_wire_2770});
or_n #(2, 0, 0) OR_589 (c6288_wire_1322, {c6288_wire_412, c6288_wire_2771});
or_n #(2, 0, 0) OR_590 (c6288_wire_1327, {c6288_wire_413, c6288_wire_2772});
or_n #(2, 0, 0) OR_591 (c6288_wire_1332, {c6288_wire_414, c6288_wire_2773});
or_n #(2, 0, 0) OR_592 (c6288_wire_1337, {c6288_wire_415, c6288_wire_2774});
or_n #(2, 0, 0) OR_593 (c6288_wire_1342, {c6288_wire_416, c6288_wire_2775});
or_n #(2, 0, 0) OR_594 (c6288_wire_1352, {c6288_wire_403, c6288_wire_2777});
or_n #(2, 0, 0) OR_595 (c6288_wire_1357, {c6288_wire_404, c6288_wire_2778});
or_n #(2, 0, 0) OR_596 (c6288_wire_1362, {c6288_wire_405, c6288_wire_2779});
or_n #(2, 0, 0) OR_597 (c6288_wire_1367, {c6288_wire_406, c6288_wire_2780});
or_n #(2, 0, 0) OR_598 (c6288_wire_1372, {c6288_wire_407, c6288_wire_2781});
or_n #(2, 0, 0) OR_599 (c6288_wire_1377, {c6288_wire_408, c6288_wire_2782});
or_n #(2, 0, 0) OR_600 (c6288_wire_1382, {c6288_wire_409, c6288_wire_2783});
or_n #(2, 0, 0) OR_601 (c6288_wire_1387, {c6288_wire_410, c6288_wire_2784});
or_n #(2, 0, 0) OR_602 (c6288_wire_1389, {c6288_wire_411, c6288_wire_2785});
or_n #(2, 0, 0) OR_603 (c6288_wire_1400, {c6288_wire_454, c6288_wire_2786});
or_n #(2, 0, 0) OR_604 (c6288_wire_1405, {c6288_wire_455, c6288_wire_2787});
or_n #(2, 0, 0) OR_605 (c6288_wire_1410, {c6288_wire_456, c6288_wire_2788});
or_n #(2, 0, 0) OR_606 (c6288_wire_1415, {c6288_wire_457, c6288_wire_2789});
or_n #(2, 0, 0) OR_607 (c6288_wire_1420, {c6288_wire_458, c6288_wire_2790});
or_n #(2, 0, 0) OR_608 (c6288_wire_1430, {c6288_wire_445, c6288_wire_2792});
or_n #(2, 0, 0) OR_609 (c6288_wire_1435, {c6288_wire_446, c6288_wire_2793});
or_n #(2, 0, 0) OR_610 (c6288_wire_1440, {c6288_wire_447, c6288_wire_2794});
or_n #(2, 0, 0) OR_611 (c6288_wire_1445, {c6288_wire_448, c6288_wire_2795});
or_n #(2, 0, 0) OR_612 (c6288_wire_1450, {c6288_wire_449, c6288_wire_2796});
or_n #(2, 0, 0) OR_613 (c6288_wire_1455, {c6288_wire_450, c6288_wire_2797});
or_n #(2, 0, 0) OR_614 (c6288_wire_1460, {c6288_wire_451, c6288_wire_2798});
or_n #(2, 0, 0) OR_615 (c6288_wire_1465, {c6288_wire_452, c6288_wire_2799});
or_n #(2, 0, 0) OR_616 (c6288_wire_1467, {c6288_wire_453, c6288_wire_2800});
or_n #(2, 0, 0) OR_617 (c6288_wire_1478, {c6288_wire_496, c6288_wire_2801});
or_n #(2, 0, 0) OR_618 (c6288_wire_1483, {c6288_wire_497, c6288_wire_2802});
or_n #(2, 0, 0) OR_619 (c6288_wire_1488, {c6288_wire_498, c6288_wire_2803});
or_n #(2, 0, 0) OR_620 (c6288_wire_1493, {c6288_wire_499, c6288_wire_2804});
or_n #(2, 0, 0) OR_621 (c6288_wire_1498, {c6288_wire_500, c6288_wire_2805});
or_n #(2, 0, 0) OR_622 (c6288_wire_1508, {c6288_wire_487, c6288_wire_2807});
or_n #(2, 0, 0) OR_623 (c6288_wire_1513, {c6288_wire_488, c6288_wire_2808});
or_n #(2, 0, 0) OR_624 (c6288_wire_1518, {c6288_wire_489, c6288_wire_2809});
or_n #(2, 0, 0) OR_625 (c6288_wire_1523, {c6288_wire_490, c6288_wire_2810});
or_n #(2, 0, 0) OR_626 (c6288_wire_1528, {c6288_wire_491, c6288_wire_2811});
or_n #(2, 0, 0) OR_627 (c6288_wire_1533, {c6288_wire_492, c6288_wire_2812});
or_n #(2, 0, 0) OR_628 (c6288_wire_1538, {c6288_wire_493, c6288_wire_2813});
or_n #(2, 0, 0) OR_629 (c6288_wire_1543, {c6288_wire_494, c6288_wire_2814});
or_n #(2, 0, 0) OR_630 (c6288_wire_1545, {c6288_wire_495, c6288_wire_2815});
or_n #(2, 0, 0) OR_631 (c6288_wire_1556, {c6288_wire_538, c6288_wire_2816});
or_n #(2, 0, 0) OR_632 (c6288_wire_1561, {c6288_wire_539, c6288_wire_2817});
or_n #(2, 0, 0) OR_633 (c6288_wire_1566, {c6288_wire_540, c6288_wire_2818});
or_n #(2, 0, 0) OR_634 (c6288_wire_1571, {c6288_wire_541, c6288_wire_2819});
or_n #(2, 0, 0) OR_635 (c6288_wire_1576, {c6288_wire_542, c6288_wire_2820});
or_n #(2, 0, 0) OR_636 (c6288_wire_1586, {c6288_wire_529, c6288_wire_2822});
or_n #(2, 0, 0) OR_637 (c6288_wire_1591, {c6288_wire_530, c6288_wire_2823});
or_n #(2, 0, 0) OR_638 (c6288_wire_1596, {c6288_wire_531, c6288_wire_2824});
or_n #(2, 0, 0) OR_639 (c6288_wire_1601, {c6288_wire_532, c6288_wire_2825});
or_n #(2, 0, 0) OR_640 (c6288_wire_1606, {c6288_wire_533, c6288_wire_2826});
or_n #(2, 0, 0) OR_641 (c6288_wire_1611, {c6288_wire_534, c6288_wire_2827});
or_n #(2, 0, 0) OR_642 (c6288_wire_1616, {c6288_wire_535, c6288_wire_2828});
or_n #(2, 0, 0) OR_643 (c6288_wire_1621, {c6288_wire_536, c6288_wire_2829});
or_n #(2, 0, 0) OR_644 (c6288_wire_1623, {c6288_wire_537, c6288_wire_2830});
or_n #(2, 0, 0) OR_645 (c6288_wire_1634, {c6288_wire_580, c6288_wire_2831});
or_n #(2, 0, 0) OR_646 (c6288_wire_1639, {c6288_wire_581, c6288_wire_2832});
or_n #(2, 0, 0) OR_647 (c6288_wire_1644, {c6288_wire_582, c6288_wire_2833});
or_n #(2, 0, 0) OR_648 (c6288_wire_1649, {c6288_wire_583, c6288_wire_2834});
or_n #(2, 0, 0) OR_649 (c6288_wire_1654, {c6288_wire_584, c6288_wire_2835});
or_n #(2, 0, 0) OR_650 (c6288_wire_1664, {c6288_wire_571, c6288_wire_2837});
or_n #(2, 0, 0) OR_651 (c6288_wire_1669, {c6288_wire_572, c6288_wire_2838});
or_n #(2, 0, 0) OR_652 (c6288_wire_1674, {c6288_wire_573, c6288_wire_2839});
or_n #(2, 0, 0) OR_653 (c6288_wire_1679, {c6288_wire_574, c6288_wire_2840});
or_n #(2, 0, 0) OR_654 (c6288_wire_1684, {c6288_wire_575, c6288_wire_2841});
or_n #(2, 0, 0) OR_655 (c6288_wire_1689, {c6288_wire_576, c6288_wire_2842});
or_n #(2, 0, 0) OR_656 (c6288_wire_1694, {c6288_wire_577, c6288_wire_2843});
or_n #(2, 0, 0) OR_657 (c6288_wire_1699, {c6288_wire_578, c6288_wire_2844});
or_n #(2, 0, 0) OR_658 (c6288_wire_1701, {c6288_wire_579, c6288_wire_2845});
or_n #(2, 0, 0) OR_659 (c6288_wire_1712, {c6288_wire_622, c6288_wire_2846});
or_n #(2, 0, 0) OR_660 (c6288_wire_1717, {c6288_wire_623, c6288_wire_2847});
or_n #(2, 0, 0) OR_661 (c6288_wire_1722, {c6288_wire_624, c6288_wire_2848});
or_n #(2, 0, 0) OR_662 (c6288_wire_1727, {c6288_wire_625, c6288_wire_2849});
or_n #(2, 0, 0) OR_663 (c6288_wire_1732, {c6288_wire_626, c6288_wire_2850});
or_n #(2, 0, 0) OR_664 (c6288_wire_1742, {c6288_wire_613, c6288_wire_2852});
or_n #(2, 0, 0) OR_665 (c6288_wire_1747, {c6288_wire_614, c6288_wire_2853});
or_n #(2, 0, 0) OR_666 (c6288_wire_1752, {c6288_wire_615, c6288_wire_2854});
or_n #(2, 0, 0) OR_667 (c6288_wire_1757, {c6288_wire_616, c6288_wire_2855});
or_n #(2, 0, 0) OR_668 (c6288_wire_1762, {c6288_wire_617, c6288_wire_2856});
or_n #(2, 0, 0) OR_669 (c6288_wire_1767, {c6288_wire_618, c6288_wire_2857});
or_n #(2, 0, 0) OR_670 (c6288_wire_1772, {c6288_wire_619, c6288_wire_2858});
or_n #(2, 0, 0) OR_671 (c6288_wire_1777, {c6288_wire_620, c6288_wire_2859});
or_n #(2, 0, 0) OR_672 (c6288_wire_1779, {c6288_wire_621, c6288_wire_2860});
or_n #(2, 0, 0) OR_673 (c6288_wire_1790, {c6288_wire_664, c6288_wire_2861});
or_n #(2, 0, 0) OR_674 (c6288_wire_1795, {c6288_wire_665, c6288_wire_2862});
or_n #(2, 0, 0) OR_675 (c6288_wire_1800, {c6288_wire_666, c6288_wire_2863});
or_n #(2, 0, 0) OR_676 (c6288_wire_1805, {c6288_wire_667, c6288_wire_2864});
or_n #(2, 0, 0) OR_677 (c6288_wire_1810, {c6288_wire_668, c6288_wire_2865});
or_n #(2, 0, 0) OR_678 (c6288_wire_1820, {c6288_wire_655, c6288_wire_2867});
or_n #(2, 0, 0) OR_679 (c6288_wire_1825, {c6288_wire_656, c6288_wire_2868});
or_n #(2, 0, 0) OR_680 (c6288_wire_1830, {c6288_wire_657, c6288_wire_2869});
or_n #(2, 0, 0) OR_681 (c6288_wire_1835, {c6288_wire_658, c6288_wire_2870});
or_n #(2, 0, 0) OR_682 (c6288_wire_1840, {c6288_wire_659, c6288_wire_2871});
or_n #(2, 0, 0) OR_683 (c6288_wire_1845, {c6288_wire_660, c6288_wire_2872});
or_n #(2, 0, 0) OR_684 (c6288_wire_1850, {c6288_wire_661, c6288_wire_2873});
or_n #(2, 0, 0) OR_685 (c6288_wire_1855, {c6288_wire_662, c6288_wire_2874});
or_n #(2, 0, 0) OR_686 (c6288_wire_1857, {c6288_wire_663, c6288_wire_2875});
or_n #(2, 0, 0) OR_687 (c6288_wire_1868, {c6288_wire_706, c6288_wire_2876});
or_n #(2, 0, 0) OR_688 (c6288_wire_1873, {c6288_wire_707, c6288_wire_2877});
or_n #(2, 0, 0) OR_689 (c6288_wire_1878, {c6288_wire_708, c6288_wire_2878});
or_n #(2, 0, 0) OR_690 (c6288_wire_1883, {c6288_wire_709, c6288_wire_2879});
or_n #(2, 0, 0) OR_691 (c6288_wire_1888, {c6288_wire_710, c6288_wire_2880});
or_n #(2, 0, 0) OR_692 (c6288_wire_1895, {c6288_wire_697, c6288_wire_2882});
or_n #(2, 0, 0) OR_693 (c6288_wire_1900, {c6288_wire_698, c6288_wire_2883});
or_n #(2, 0, 0) OR_694 (c6288_wire_1905, {c6288_wire_699, c6288_wire_2884});
or_n #(2, 0, 0) OR_695 (c6288_wire_1910, {c6288_wire_700, c6288_wire_2885});
or_n #(2, 0, 0) OR_696 (c6288_wire_1915, {c6288_wire_701, c6288_wire_2886});
or_n #(2, 0, 0) OR_697 (c6288_wire_1920, {c6288_wire_702, c6288_wire_2887});
or_n #(2, 0, 0) OR_698 (c6288_wire_1925, {c6288_wire_703, c6288_wire_2888});
or_n #(2, 0, 0) OR_699 (c6288_wire_1930, {c6288_wire_704, c6288_wire_2889});
or_n #(2, 0, 0) OR_700 (c6288_wire_1932, {c6288_wire_705, c6288_wire_2890});
bufg #(0, 0) BUF_1 (c6288_wire_32, in1_net_0);
bufg #(0, 0) BUF_2 (c6288_wire_57, in103_net_0);
bufg #(0, 0) BUF_3 (c6288_wire_62, in120_net_0);
bufg #(0, 0) BUF_4 (c6288_wire_67, in137_net_0);
bufg #(0, 0) BUF_5 (c6288_wire_5, in154_net_0);
bufg #(0, 0) BUF_6 (c6288_wire_2, in171_net_0);
bufg #(0, 0) BUF_7 (c6288_wire_30, in18_net_0);
bufg #(0, 0) BUF_8 (c6288_wire_10, in188_net_0);
bufg #(0, 0) BUF_9 (c6288_wire_15, in205_net_0);
bufg #(0, 0) BUF_10 (c6288_wire_20, in222_net_0);
bufg #(0, 0) BUF_11 (c6288_wire_25, in239_net_0);
bufg #(0, 0) BUF_12 (c6288_wire_330, in256_net_0);
bufg #(0, 0) BUF_13 (c6288_wire_3, in273_net_0);
bufg #(0, 0) BUF_14 (c6288_wire_6, in290_net_0);
bufg #(0, 0) BUF_15 (c6288_wire_78, in307_net_0);
bufg #(0, 0) BUF_16 (c6288_wire_81, in324_net_0);
bufg #(0, 0) BUF_17 (c6288_wire_84, in341_net_0);
bufg #(0, 0) BUF_18 (c6288_wire_37, in35_net_0);
bufg #(0, 0) BUF_19 (c6288_wire_87, in358_net_0);
bufg #(0, 0) BUF_20 (c6288_wire_90, in375_net_0);
bufg #(0, 0) BUF_21 (c6288_wire_93, in392_net_0);
bufg #(0, 0) BUF_22 (c6288_wire_96, in409_net_0);
bufg #(0, 0) BUF_23 (c6288_wire_99, in426_net_0);
bufg #(0, 0) BUF_24 (c6288_wire_102, in443_net_0);
bufg #(0, 0) BUF_25 (c6288_wire_105, in460_net_0);
bufg #(0, 0) BUF_26 (c6288_wire_108, in477_net_0);
bufg #(0, 0) BUF_27 (c6288_wire_111, in494_net_0);
bufg #(0, 0) BUF_28 (c6288_wire_114, in511_net_0);
bufg #(0, 0) BUF_29 (c6288_wire_42, in52_net_0);
bufg #(0, 0) BUF_30 (c6288_wire_117, in528_net_0);
bufg #(0, 0) BUF_31 (c6288_wire_47, in69_net_0);
bufg #(0, 0) BUF_32 (c6288_wire_52, in86_net_0);
bufg #(0, 0) BUF_33 (out1581_net_0, c6288_wire_1955);
bufg #(0, 0) BUF_34 (out1901_net_0, c6288_wire_1977);
bufg #(0, 0) BUF_35 (out2223_net_0, c6288_wire_1982);
bufg #(0, 0) BUF_36 (out2548_net_0, c6288_wire_1985);
bufg #(0, 0) BUF_37 (out2877_net_0, c6288_wire_1988);
bufg #(0, 0) BUF_38 (out3211_net_0, c6288_wire_1991);
bufg #(0, 0) BUF_39 (out3552_net_0, c6288_wire_1994);
bufg #(0, 0) BUF_40 (out3895_net_0, c6288_wire_1997);
bufg #(0, 0) BUF_41 (out4241_net_0, c6288_wire_2000);
bufg #(0, 0) BUF_42 (out4591_net_0, c6288_wire_1933);
bufg #(0, 0) BUF_43 (out4946_net_0, c6288_wire_1936);
bufg #(0, 0) BUF_44 (out5308_net_0, c6288_wire_1939);
bufg #(0, 0) BUF_45 (out545_net_0, c6288_wire_75);
bufg #(0, 0) BUF_46 (out5672_net_0, c6288_wire_1942);
bufg #(0, 0) BUF_47 (out5971_net_0, c6288_wire_1945);
bufg #(0, 0) BUF_48 (out6123_net_0, c6288_wire_1948);
bufg #(0, 0) BUF_49 (out6150_net_0, c6288_wire_775);
bufg #(0, 0) BUF_50 (out6160_net_0, c6288_wire_781);
bufg #(0, 0) BUF_51 (out6170_net_0, c6288_wire_1951);
bufg #(0, 0) BUF_52 (out6180_net_0, c6288_wire_1953);
bufg #(0, 0) BUF_53 (out6190_net_0, c6288_wire_1957);
bufg #(0, 0) BUF_54 (out6200_net_0, c6288_wire_1959);
bufg #(0, 0) BUF_55 (out6210_net_0, c6288_wire_1961);
bufg #(0, 0) BUF_56 (out6220_net_0, c6288_wire_1963);
bufg #(0, 0) BUF_57 (out6230_net_0, c6288_wire_1965);
bufg #(0, 0) BUF_58 (out6240_net_0, c6288_wire_1967);
bufg #(0, 0) BUF_59 (out6250_net_0, c6288_wire_1969);
bufg #(0, 0) BUF_60 (out6260_net_0, c6288_wire_1971);
bufg #(0, 0) BUF_61 (out6270_net_0, c6288_wire_1973);
bufg #(0, 0) BUF_62 (out6280_net_0, c6288_wire_1975);
bufg #(0, 0) BUF_63 (out6287_net_0, c6288_wire_1185);
bufg #(0, 0) BUF_64 (out6288_net_0, c6288_wire_1980);

endmodule

